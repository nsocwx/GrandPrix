PK    S�U&!S  �     cirkitFile.json�]K�۸�+[�UT�rn����vզv�
$�V4�D�ػq���^_j�!�V�s�g��l|�@}���g��g�����M�ZN��N��:�b�����\Ϋ����yy�<|�G�/6�V�/��]Vsm
b�I�"FQ��2�I��il�xN&��P�h%Ef#Q�$2&Qn��L�=��Oӫg���ff�fF���(ir)�37��(����̲"�x�c\`f昙%Nd
7\�Ǹ�	n8%��9	wʑ�r�B=�)�@Y	]���DEF�d"���p��
35�:"1Oc��(֑
Ð
Ð
Ð
ÆD*2'z�"�K'�8f�I��Lf��JfsJ�C�L��5���i��i��	]��.ǆ6H[ϑ������C�,�U C����A8bf��y�G�f�1��P�<��fZ�̐,׹�X��H�L,Y�<MK��\g`��*t��w\a�� fJ�@��y��k�m:���Dq��(��I�� :�2MS��,�|`0���/1�!A�=� ���!�F�K�0>r�m��5�:Q&h��Ԑ����!�:��@3��@ˍ�{�j��j�Z#k���$���b܉�B��Ɖ��J��
j*��	����Bs��*2�� Tt*q*I*��!CÐ	_�Ða����q�c�l!�g�0d�`�� N$!�M�0(faP� ��(V&f*Ð	�b��0���A1c�Y�0(�aP��al1�b~����E����Fh]p<n���Ɲ�^�ɀł��<���/��6�B�Z�1,�F5�,�%�q�B�?gVX�9����ȸA�g�,<�?��0�]hA`��Cs�q����҅��8�ޛ�T�z/�k�6dꍧP�A�� Td**�J�Ju���4|i��0 �aL�@���0b�,�Y �,�Y�0(faP� ��A1�b�<�y�P"�y�(��x*g�	�z㩜]%pꍧrV.��O%�\΂�z㩜�.4��S9/]hꍧrV.��{�
8��S9�D��O���.�^�߫�����<P=�|)�v3Y�q�ܥ�unד��ןJ��b�?@���t���XG����sR��z�D���*5�s�z s�c�o��гB�Oo�`�bB�[`z��Kb��a�[@�co�X�Pc`j`����`�z@�p�ڢ�������|5 s�����^z84�yZL�����:�}�HpP�p����t�L$��?��}^}v��Y�}9�G���%����C�#e�i!�lv�� �(���(w��9�C�2��!
��d ��$�dZy;�˚�����1�G�;����۩4��)��b��%V��,�9M�C*�!D��	�`tC��7�8*�!�U�7� �;TkF$p��wx����qN�E�A8 ���a�L�%D�%@V߸Zp.8�K]i
��3�1B��n蒂��Ri��V��_�������UQLb^�{���`���K��Ls�՘;��Ut����2��S��9>F�O����0(K �������PS���7_Z�P����KKk\��!��-�aa˺����bX3�-eXcʰ8eXsʰ��X`r,09��c�)�"�� |]f���V`�,��d�9�w�a��0o��nO������$��K��F^�z#�՘wC���젗e`�5�
�����0���yX�^ՈC_��hշ��H��}��o|�1�=�^D^<�|��?�WW��+��U�eY�J�H��R߹�S��2��S?��̏`5m?��̏`~�#����Gp?�.<�?���ߘ�@A���@��ꗅ���Y*u�@�f;�u������Hc;ّ4qR��"R��q,2���+�i��R��?�x�*�#�(�ͨ\�BD%ʺO�H�9�+�s⤜(���R��)(�L���^(��q�z*�K��/�H��i�ua��.�뮉�"e*�i:x�Bi+���v|KYP����ՍtP/��]��Z��o}�˱�=�:����_�W��nu}2��ԸK5]����䍓n�zc8&Ý��F����]8���7���{l�t�g�q��}��S����I����l|����~�rk5�]�6�]��6�]��6Ż��۔욒NS]ٯ9$�ajצ�Mzפ���}h�h����Y,��ښ<]����P��rSyP�B�Dk4a��F�_Y�B+g�,t������~��?>_آ�#�~������2�G֫��J['�/K����vS���o�I�����[���f�����nQ���d�~�<���_�st'�Yl�k���/�L������\[�V��4���0Y����1���l�,p�_�ڔU�5�#�gr�5���Jr'M����O�R.-�I�D$�����sB�>"�t�We��v(��NV��-��23y}qe�:[��~�(a�A�ȧ��-$�N-�5[x�E6[T�%&�Si�%r�M��q.n#���8�;�)�����jʩ)����Bj�hDD#Ј|F�3"�a�ZB�T�����k���m�w�������.���׼\�����	��qv��H�t�=U��D.o�?T&��M�	S�)������2iM��J�"cGF�8R2�N}�������DcY��d���x��ڄ��fS��L�<m��r���T8�r��;)7*���e���q�]���8�g�7q�(���Tz��6Iܿ�6�ͭS��@�HX	�&ܧx�q�vN�/nC�Y�'BI�q���NE�=�q1��EG�j@�L쬖�����md�	�}����:D^�P^�<
�M�~-�~\�~�{����R����[O��3AO�j��S�p��D��Hc"���b����j���	�L@"�`��k_�(�{#�Xy�^ZʩvJ��ESi�Y�&��[�LM��N&��4-t�ٶ@�V�y���5�����E(�Yٝ7"r'[ȝ�:��u��4qf��G�<�$�Qb
�����u8A ���F@����`�n!P+e;G�S��{'�o�����}~��П�#k��q\�_Me�?��>���b4/��Y��⇏������t�M'Ţ|y��d?�ٯe���0w=�q���߿�W�����K�vL�i�9>�_��g����߿�����&��:LCG����0����[|�s]�����m/�C�('g�Rj��n���d��O��{m%�3�(��t��Oc-gT�N�t���(T�L�ԩ)O�(�����y�\n׊���� �]���ݴ�ݪ\|���zxO=�|�IHL�r)�ӻd�c=#�Ƃ�.��"��!h3�O���}������j(��m��yN�\�O�T��[+]rU�VA5�DZ���Z����^�������-���Ɍ)�U�	I��j*(��Xk�e�9cB��"�@ԟH#r+�)W���xGedD͸"���K�US��L'��XM]�*��:q�WE���1P�`�r�D����,G���w���x[���%�Փ'�~�_�'[���:���U����q:�?3l�'���p����V����˯����|���I���������B'�Gg!�ک��Ǽn��TdM�.�QR�Ù5����sH�����eU:e�������ǉ?����~�����������>�0��N�q����n��l����n\�+���L�ӭް��������)Զ_'j4�X`�ѠPcA��e?�N�Qݿ���n럴��N��_<
��3C�S�p]� Cpw!�N�<�Z��V/����to�M����;��&и��7�F�np2`^�5�䀱j�����w	�4/1$����`(�X���\���<-�&a�"���	�.��M1T��<.Ԡ}9�����:�4'Y"6x`l����A\Ȣ�k���+�=�nC��S	�U8p\��_�Z(p\��ק������A��)zM��S��n�ٱn�PS&f*i�,΁��l�8й�=�����(yE������N�!+	�ː0+�	G��A����Q��>.��e��b�z��F9���]���\ﱗ쉒���d�]�}3����|(��}�R'������A���6���= ����Ft`�!8w�bH0�N{q��*rE/����&��R�,h�`��C��+0���ႛ�}��`�x�F`�/�D���2��0do����2m�^ы���`������ʚ,g��A�gXB�ov��2,W�o {���jX.Z�$İ�F������!�_�+��(�F�o �m[����*���?�-��,6��M�G�_���,_��o��+��y�_�6��?PK   �jgUD�#��9 �9 /   images/44ae2a6d-294a-417e-8c08-7c32f15c3a8c.pngl�eP\A�-:�����w',��3�%����w�<�27�[���N��ǮU���cW�Z�O���<*)*  �PT�� 
  8] �+�0� �%/��"?��@�y�� hHD{1G���(� �����F��- X���{���(R��=����ތ�����J�1�%�y�+���@fT��F����x��ۭ��q�gu?���F�s�>��Y��l��d���ZG̦e;���g�����hy��D[M/�{wm�㩮���]OɄ�o�LW#m�g]�ț�5ܛ��S�Ż��\���H�߸d����'�����լ�t��
����$�)<��PJ *ڱ�tô�#�=���h�a��s�a���i��b�P�o�y��j�1��!Zn&9���|�v���k3K�|�^'�_UiGri����;'܏��4՜�I�<�r�Po_����/!k���Gp����vs	c��Pѥ�@�{w�����>�e�-����j�s��:�-�p0�m�.b�
VNl@=�6ک�A������v(� �/�s�ʕ	hn�خ��v-'v��''��v{>�z�u$�j�.F�h�ulr�aX~�;�QQ8H��g�(G�1���i!L��*N^%.����^2#>���Q�FZ����I�uQ�'�*��w�g�&N��+TU��C����g؃8��a�,܄�|op
.z%^鲍.Cȇ��ja�<��M��T��n]�\˻������RQcF�E�ϕn�������e�\X�"�A#1{�������:]B]\顴���
jע�����e$l���a)��d�L%'� �Pt����1�	�e�0�#�P-�&��i�n����7��*(�U6���3��C?&7�_���eM�~	l�I�ŭ�@��C�Ɉ_rg�d��s��zQ�&��R{+�����h���/�kς��W�^O�����	H�N�>��
�����5�+�ԋ�-I��.Ɏ/C���ET%妕�h��h`�4�JC����_�Sp}�����TJ�/�mI�H@��is6.��.�{d}6-��E����s�*&a�OLb��ۀ̇_L�x�0�Ԁe�U��g'@M�q!G� �{~���; �j���+��Gŝ톩�Ƕ�Q>��laG���.�64�1p����/��^����Ѕ�J"�P�Y:��|���͐�9	�Nx�N�(ԀaӲ+�8�A��N��+q���$�U���Z7ʱ��"���E���[`#�A;����P�d�G�v�8��ت��Φ �����u!���'��~��(ޮ���9
?Rnݾt:i�;J���lv��Xc�2jW��T��D/5����>�KB��!v��M ˬ��1��5,���[���� FvEI�	��a΅T/�Ra�\��)�5lO��N�������!es��EC�� ~�B�l��������߁��e H��B�'�j]��Ce֐/���V�k��p>�G��q�bW��N!�?����
� ּ��@8B�.��6ʆ��<J,G�D�����s�d����'J��P�E	��x�x9�Ô�l
|��_}��3u�����8�\|;+O��%��V���V�ݩ��M�n�]�_�
[Vݺ��X��ĸ�w���u
3�!��a��-�MZA�o��,Ii'mF%LB���`j$*0gU�YE�4m+5t"��Rp�T�*@Q�pkSQ|��,xFe�7���~W��g��ӊ_`���x��	 �n%�]�2�C t��p�Tp�T�(�s_�Ҹ�~�5��"]�"Em���)�0f��MQȓ��vfS�e���q��e�:�?+ Da�Z!��i[�}S~IC#�U�i2uM�;�L�A�6Sw��;�d�6@���tz�Ѻ�E�?L|�C �$�Q��;�?��X@��2y����#��3�;2G����P�ۣ������yܾR�?W��zbVʼ�m0��A�Hʬ���-��x��?�O#5!s�|�lVt�b���W�3����0l�11K�g�_ʕ����Ӱ�$��J��HQ���H��f����e5f����s�^J���?u�2��_���|����r��W�� ���S%�l��3��S+��$��5_��(ע9�p4��{K!��Ɵ�r��%��_��*�ܳ>������](a=����Clj�N���~7l�}uC�:LUJ}O�@]g�$������R�x�4��`�e��uuռ3�����s�Ƚ;l/��6��#������xB^$(�K��:�����!�
_'>���7���/�3�hHSssr�^�J\cP�48�԰�A�EZ6��Z��lr��a��aք�9sI��'�ռ5;.p�F�UAsNҶv�h�V'}�}��!�H_U���hF�d�H���_��w�`��w*���B�9{NN��i+u���"%�Io��b9�hE-B;���R��x}��9�@��R,E7�
 ���\'�*1C(�gϟ|��4-�_��;r(:�*�Q��k�]P3'K��-ݪH�i��U���\g�ŦK��ؗ���/R�@���4d��г��o��\L����n�}nB�k���<�͛Ωo��6Q�C����E���GKUd~w��6��Vu(i�X��Nuy���u=*�~3����A����~�6���ӗ�3Ζ��K'�8)(�M��U��)#����L;�h��/���6�lx��㨺��<��A"��L)����$�� J!�%�&�#C�f��~��yJ�x�벮n5f*���}�ۯ��?'d�w��W7�Gz���/��^S�v�p�ض4B��R�F��c�>��"J$� ����^m'!�������,���
�+mcŦҀ�f��'�����܋�� "��ezC4�nL�ݾ-�5��Aݎ���{2Mm�4���'�4�t>0w{-�i��qg��go��~	���S2�S���|I��aT6^{�DR�8�o-�I�*��m����f�O�#E@�&[a�����oU�eRNUR�F7�/����k#���n<y}�����$Zw�k�"�3��	�I
����Z&�+Qz��Ij�r��r��3Q�ԫ�p��L֥t��(�I[͕��-Ueee����@��/�w��K�L��\2c@���Ӹ�ᩄp��)@�vÜ�;�
}��_+����;�j[o.Yw�1j��ĨX�T����Or�Z% U㧘�E��P�[{��Kl<�܅�F���A��߇�4}q󍘧9�!r�
�sz��m�ٜ�Q����~����w������ۜɭ}� �ѥ��X�~@��2o��t�X�{����B��:qQ�!M<�N)p&��hRt�r�a8���?3���R�\��������a�a�f�H[	;�ҬHwz�G�8V�_��<}�`V�^�u�!P�cV�[1�Yn=��U�"�/�3=H�:fI��/�Q�+a;@�?3������C�1�q2����}���He$�t��܍wU�<G=#Di�#�hQ��=дP�\�<��5������H�n�M�N��Q%>l�^�{^���9���	>��Om����?X"�$��P�2o�ג��(kr�eG���R�.-4AKlM��!otBj)���~�'�n� ��`<�y���e�5Dɘ��B�((W��FVT;QC���։v�VND�0��'\�؄t�}T�LB:�P7.8��c��>��	?�lCu�f[ 8�t�����2�5*�#d��U���*ݷCZe��EpF� ÌCAC`$_���h���}�-��˴�2�eB���B��.�.w$�d-��m9���8!';O�@�;J�L!$m�8����u0���pț�k���V��BV?�]�V�E���zR�ށE�<�C�{�{#&l��mz�g��) ��yG4�PiI�5�H\���#�菭�͙`,t�y,0֗�c���<�MᏙb����H��)���|�Di�qti��h�ػ[���S��J�6<��YaB<i$)4��S�g�#���iI��p�����0Cϙ�����H�9n�uh�#��?�P���]'�*:�q�0&iŴo�Q��������&�2�l hv,���	�kP����͝|7}8�n��H�Í*zm1�T���`i��S~H����=]m�+���x����ID�vɊw!n��Gj�!�K-�jܺ{)�n����5��F ;�<>�z	��yw'���N�i�ؼ������C�FtJ=��;)�+TÌ	��we��g�u�Z3$�8�+sa��^K�f�pm,d��h!�>��7	���YpTTTHL��X���q�#�t��!m!��dg;�r�X��?Mё�����k��>�����m�@�f~]D/)� �c{�0�P������@�j�x�sf>�_������5B!J���x������ֻ���+0RS����{�P��Y�8�k��Y�����*��m�Rq3瑅`P��[8@��oɬL���d�L��w���:�E�vq��@�ZSaS�O�{�����t.�Z�K�N5ʞ��n؄��,��N=%��g�R��ȄIDb�L̽/"�֒��㌃�V�]�o���BR�g����/.1�-7	������I{G��%�$�,Ge�����T�؊��V�:r�'`3���&� �c��!�fʂ����5GoI�IWMM:�)~�;����+���F�g�z�I���z�
{�e?�Ck�����d�f��r���r`)��s3a�&���?	���Q%�$F�ߖ��%��n�K$�R���!��g�n@��L�i�L��xаN��D36�_����%nF>$Up����@��Ǡc�C���U�m)��M�:���HPH5_3K�Z�Ɇfg�N;F�n��Nc�U[��k'�VC'����JY�5Y!9g��B�'�ٗ�lY����>�{����	Z�p� k)$��q�OYp5�1�k����*t=��1�/�#�$`5�-�c-�$���2�>sGk���#QI�-���#T9�K��ɭZ�@�6k������iX$ٿS�@�1��;6yn7���U�|��t��;r��q�������,�#�'����a���������?�gz��w�ay5��Z�������!G��\p�����wo�~?z(_�6J�Y[�S��n�{��Kx��n��ϟ�?`�=��R-`��3����B�R$�L���Q7�L�B�N]�K�?�Q�!��?Xr$��R'����N��l�B���������LuZx"�$�B��s"�Q��t�6�aw�j�!_��[\��bVz=�!��p��T]�2 Օ�uA�k���3Ȼ�	�=$�#'��a�t�G��"�"f��Be�a��[�1+ܖzeojIf�o��=���T�I�c�Ļ/'W�Y=��4�>����du$����s��Q��&�M��7�a�B,5�E��}�#�l^���gMep�i��A��pjq����|�zU��f,r��j�q������6�R��޴�݉���0��m���N�!���X��Wg>Y�;�Q����������CQ��X�F��+� �Y0�Ra5]�l���������=�N����M���Q��4�9B��Y��wkqP>��<D��ٖ���$`m�{K�0��E�O�?4u!�9AY�����o.8V�Of���xHN<d�Ӱ�N��4j�T�o�Mk�mk(���1��³��A�.CU��x�������!����b�W���H/X�B�F�X�k��y�^p�ҹ�܋��>/������@�F�W�����򿓝�C��#�>{�}6�X+#�����{%�{%�Ö{��T�l�Є3ӘA�����Cwęg��Q�
��?�K�Ӓ�w�<|ځ�;��"��V��A��[�U��^�U��Ǿf�-���RJY��LF��6g �m '3pRݨ�������;��Do$��	���s�����S�K���V\�7�����n%�^�&dF2�H��� �p���o��N;	6#
��U>z���� ���V�`��m�y��ۿ�dD���Iƭx�#��~��ܭx�����Qg׿s+m�Ț�g���hEshKx�{b&Ȼ/�����C~��ԟ�T#*ثɓ�kY+"�� ':�$>���$��`�qV*�|���P0��!Q\`oU�	�
iJ�V�j��&��n٢�Ә�c�/OBp�D֧�X��:��󓴙���co�
���/�������H�)��:Sr16����	���e
;y��R� �� 4�������K�8����1��G�xXt2�v�U��@+V�������)ӂ"�-Q�>j�#���G�ɠ�,���| ������7�)�����z��s�e]�u�X��=���^+3u���ĤW�$� �a�_j��ɪdWb�}N)��#I���x����ZASJvds���)3&$ɀ�_�]�n�D4&�P��i�X�����4VQ\��h���ӈH@Q&�TZɂ��G����<��Pf��4l;��U���iR��~_� ��}bllc���Z�����뾠��Y3||~_.A�_|��_|.|��h#�� �!�	N'o�#L�����j�
��x,��P��RpB�r������h֚�ɬ��br��-1&k�Ms��)�<m�{�� �7yZ�7_*s����B0B]�Z��`X������j�2����f����yo�,��N����P���v?:�u�����0�'=�.>U���gn���@�J�r�z8�^����c��!|ǅ��E]鋩s#M{�ʑO0��8$�=Ėw/�����e���M��n�_������W��G�S��:�����"{����w-���Y�#�1�|o@�ݾ|k@}�N7���7u����n��.�� rS�]n�&�N��]��̤�#|F�4�9U���@�����&��,O�
eG���1% ]���b@*��~�g X�k��_9仏F��z��M|{|V�y��3p���#����!��W"ʣ�|��|P�&�@|��[)���G6�����pn�[`�0z��w���:mw�D� ����`�9�D8Ұ��g$H���[$�2�9Û��x���`u�n/���0s�{0��������W�c�L����'S�u�}=�U�1��ۤD�M�5��c�Ga^�Ӥ �I{�5L��巄<�A��7W��2v�����L�z�Ȳ�yR��A�N��GD
�;�S���t�Q��J�%�#�oހ�r�1AV���&���W�A�:�;~g��jT��(��d�H�Lt&|ӎ��i�d��~��pl��?��s�cNХ�����exE?R[�PԖ<�7�	��^��t��q�)�/�Z��w�_b�(��tt~F�p��"X��,��U2�&-�D1z�G-�%���zT��N{�1~4�c�d���e)f]�\���4CԳv������+��e��e�i�p[�9�Ӳ�Y�������K:}�vL��je V.
\�<4�<Ռ��tT�rf�Rj��{�#�S��6'�4?���H��I]ϋ�QOĥz�A��D�	B�`-~R��ft��� ���t��M����P��1"E��X��E�sA�Z���aI.�q�)�u#)��8�Fr-D��|&xT�D0�j�x>:�Gĝb�&����xH(�d =�G��Lл��Sk���K�b�,��|a�$��]�$ciD=���ԏ��3����ޥ��F�kvț$���?�L�9����2?f�?c�7K1|��~�r�eM�b������t���~�g�0�-	u��m�ɑ���R�(%m���������)���YB���E���H��6��FD�>�;T�_�g�����	U��K���KM�M��ҟ63��Ə�l�.V�g��p3-m���&j�s��f/���/=@�LB������*��z���aM"iSdB������bί�^���l��G^/R�؜�E �� �Ƃs:��j��~��	�p:�/+V�r�jgX�0I&S�=���*�ǐ0����좖?->DN_���u�a7�3V�R��_ɣn�����c��Z�t���n�6o:5K#T֐�����W�����
8�0�P�>�Ea��kği?i[��4��#�C7���">�"I�=X��Om�y��^Gl,@��V���w��#�qW3tc�aqud�&�o�x�6?f��WC��h�Ep�s
N4���g���d���jYpͯ����@�q�� �O���t
`�*����R#7�9�%u*y�'�W|�(w�ǌ�]�,8���e=>�� 1�UF|r���p��~�G��vo;�QpG��	�ա@�%m�����#���W3����|2ă��r�<!�I�����Uhx2�9ط*i?��,}������@%�w���-�gf|��v6�ey��\�8����/��XUY��^s:�d|���	R��g�w�oIW�ġ���4��|�	��A>��h�Qc�?���яCiR"���}��g��F��>�'��	��v����&S���B�Y�o:�yoڳ͘���ú��'� �^V����su��ڕ��1wi�?� ��0?P�%ֆ�ߠ�(Y�b����Hc�^{��AV=&��^I�l�;��W�>?qFU�~Q9��ODe��������ҙ]�x�0i��Sv�=�y	Qw=�W�N��1;l�(T�Z����ak�@�N\du�����Ɔ~�.CN�<�h�]g[E���������#����^���~����F(�ω�������k�i�����\�$���fL4�)'�a�/��Ͱ��K�[5q֡��6	��|i�I'�����%-� �f��;CR�#}�9�ʍ���?��z�~cR��<���!tm��p�hNl�o�pW[2p�qd�^x�+>������'5�V�!����>��e�N������(k|�0<_�_'I8���u/�c($���xbe �3z�Ľ�D�����nڛw�\E�|�P�qK#�l~Y�C�݄O	qœ�(�WPY�y��N��Q͘��t�WT����8�[3!GR��[s'[De�4����I���L�<�NٱJ�+��D�`�'I��:
��0W�?o?���\4�>��7��T K���F�K��#ξG�u7����B*�lS|S�y+����?N@m"�K%���RW�'F8��>}"��Bԫ��9�,�u�8��j7��׆�M@�Ñ����%@�jo�6Ri?/��<1sr����,ε�� R��4 i-`�n%o�UJ�^x��\��6�(͇&C�D�6���E�����F���)D?�o��F�O놏�e&������xZm�{���٣>� �s�\j�?��.��ޏ<׽�*��5��nG�o�a��ssa����"d9��o�F6�o6�U�6�l���ۏ�9:�U��%�ki���X�����P؊���'g��vY��e�y��^I�%V��va��9��[�@3�:��*�ܿrϵc��3�~�QX_�����ƚ��8s��3�4�0�S��}g��Ʉ�`�����Q��_���ޖ��m�7�ê!�b%73�ɐ�)��ؾK�T�*�7QV��'a��	gwh2G<�׮��_�O����@���AUj��i�d�Q�;-_ǅ��@�w�3�s� �Qs�N[8vV����/�)j3k\v�|����R��M͓-��͖�D���?��R�����e�/�m�������r`t�SuVa�ZJ��)hM��������~�I\�%�R\�dU�� Q�u9#��b��'�����Qgp(y��!��:Õ3�NcQC�e���'}��Ih� �9=;����_7C'gd����8AC�Q[�NA����������8GL��_ŹP(IW��Q��$}��vz�ԽW��g���=˰��HA��dG�l$�'ش�����1Xf�I���B,�"*J5W �M��x`�9��!g�[`j�ө#ո�wVqy�/��h��-L��qt5���:�[oy�&�t{�s�Jty	f3�������	�%�
�#���;�7�v��ބF���P���� 7;`Y��Ru�7�-7 GF�#L6�����9b4��~4s����B���p�(
�(�b��x�=T[D����>O�mOWީ~$�bhJ�W��|%�`%!�ޮ
� ^�<�M��q�d�:���$7z�Y�h��g5�ǿ�!6����	�t˿��2�,6캈{Q�R�vJrO/�Ɛ���7�C2��O��n�J�Ļ(m!^�AJ�̕��LD���!�˛�q�?֌���`ѽ-ʹw5|<u�E�>�$h�ί�I)���v~s��v�H$x![X}z�ְq|���_܏��	���s�����{�X95��>�Nٵg���L}f
�j�9���6�m�̫eפ���f^O��D�n��ܷq���P��-̎å�FES�O�Z��g/�UMۤ����ڰR��ޭ%��c5X��F�B��D��N����O��=[{�[�W�D�mX�a�> �H�"��.1L^��M����	��2����Zt�I!�"�7֞��6h��wFZQ�+#lC�/��.���ʴ8rG�\�z�߸v�X�epqs�h��	�l>����/᥼�ϏgYYL�p|����x�S�F����\i��a\�V���8"{�>aU�i�K�A-_�X����6��/Y��㲼�^���̪VIoJx���
�}N�:kc��;ц׊�����T�l9A�&�����W���7��+Dx?G~i�P~?d�Q��j"QCz�݋����i�$G��,ݕ(~�`��yI��V��G}Ho�]2]?bϗ��	�#K?�ͩ��>.<"lL��S���'R����ɻ����(!((w:'m�~Xg�ot����O[������QJ#�yB�Zo�C��X��U���ȴ�V'B0
�P��,"������5�W>N$�����+4ki�~V��5
N��N�wР����[3r/�6O�W�8�[����1�����k�|�@'����lB�e�;��)���[Qf��6���ni¼��f)��ӵ��p���n��-ސ�Ĩ��_��v�F�R/b2�(j�r�@�bz[��P$iQ8�p1<% �%�~o��}V@��z̲�h+��u����)��������#> �FJ��A �K�ױ�zpG�� �O(���1
9�NC��$�&�5�|�q��8v�5�fn(ר��y��My?���*j[�HN��M���z������#E�C<ul��2���#�jkQ�K`�5��"'�~�Փ�:�)��r��^I�H5�v;W��WT�?_(��86F�þ�y.m�.Su�f-dz�t+S�b�RY���&�r�e�̓���Sщ*���/��?g�^�OK6�-QVB�%����^`D��O˦�x��`X�K�#����ʹ�|��YK\�N�+�g����4��V������ I��V���n7xy5�߷%���1�w'�F�4�#g�b���"��:D̈���d-�6����)����f�_E�(�\�:FU�|0{�L���oX�"H���#F� *p��:֢V|�z��!e�r�����JGq5�Q��x�z^�lv��CيMՊ�!9�L�$��[
0u��<:�9[���9��KGf���7&�����j��[�-Au�Vn�/ ��_<&�G�Bۆee�?��L�$��A��X�[F�ИJM˕;��@�5N����+���<���1�h�}�����(��?����C�'���G-�S�Ӭ"�<�\4�d��jn^e��G@��������6F'}GL7���6�-�2?Q�$1�a^)��S��w�m&C#����UU̔�}�%�+5��Y��?t,����nH�Ƚ�E���>���6u��i���������j9g�kO4�*zR����	2�@P�Ɏ�3�#4��&�YY���H��oi����A�!�~���}�꾔ʧ<�je����d5�r��殳P�Y,J"��l&�'Ӯ��Ƒfed n��������y�|�b�/�D��E� ���Z�`��7�`*���ZܨP�Zn5`.-b���r��<�N�i<��R�R�v=�fAt��I�`[Xp��7��̈X�C�fC�f,q���eɸM,��z�Uu�x><�Xa��~�-�X4��h�΍�%|ݮ��Y0��?�n~KP��-�Iq��,�Ҽ=�[�F�l�y�/NX��Wt��5݄1���V��o�޼*8���Ƨv��ׇ>βZA���n6�s���:��E�E�`�?���y�d��v�԰<���!x#�28���0��͙jy5��Y_�mM��_�:L4���� {P��13�7%��T�Q������T�'?l���x&߱��f�����z���t�.�e�����s!�VN�	�e���/t�XY�._A@�R�R�K��r�o1!����1�D����r8HZ``=�� �Ӥ�C��J\|��mk�b`���L�w�/H"Y��1��Rّ8�t�e��8�,x��E����
N�B�A�[��])o�a�gj�)߿�4��P-�z�Y�oj4��V)�?��_k�KےE�B*I4�S�[�_UVr +��|9�E8���l2�!�-��iD8����a�p�Ӻ_r��wu~��ЎXp6����kWaZW���ӏ��F��J���1���D���'�}��'�5�):�i��|�~+��)���g�$���H��i����� &9���MX*�iN�l�aV[���`,]*QM����������Cm9�3st}�;k�X�8G���k�!}s�>4[�*A�b}K���=�%T�=б�c�`�y�.���wc7}a>X���#��c5�b�qoiLL�m�Q��:ofk1���[Q��_�(�쮬G!���p$#�}���f�eZk�ƺ������X��z�D�ُe�9 ��
��h>�d?ab/��a�:���OI�/�`*�.{9�A�b�2l�8����@ԗ��l�Q�+�ג��!�z���A��O������ߪ=�1�C2���a#��~�B��_���'���~����ҕĝ��M�MyJ���O؛�s������������a;g��F�׎mU��,��ޮsơ�5��[z���|W9��b�,���P��)r�,)�,�y�}(D���7�v�f��Z�_� ��Ϗ�E��ݫ��$\���	M���J�$��=T�3����S�weO�����V����W����a�%wQ�;��0��%0پ�����D�`�g��������q��K)�KF����ۓ�~�q��6����K+�萪��,ȱ��^}��R};8���^��� �{o7�����R�i��R�g�c�6�lF�b� �?<���\#</��0����M,�ߧ�C��ѭN�?���Z����\u�K��U���i�t#Q��'nR��惭��W[M��zߠWh�#��ωW�;��&#���;3��;W ?d>�*_���},}���86"G��m惏L[/�I�l��q�=�r�l7��E�I�W�)�0x",B�,���bّXebiq����Wg/����7rۘ����؏7Y�m�~��V���L�g>�O4�G./���9:q��T�m�lb�Ԋ���| ���*�qt�+��7��;�=�ldɼ��K�}�ϖ��q濆D}<��Y�g��+�&̙�BXNb2Q[��h�`�e�k� �yM�F��ĞY�\�N�����"��R��F�b ��N�;�؞cWÕ9W��V��M�s��s~9d�i��}!�����q��E�5�(�5H\3;�'������;��2Y��T8�·7P:�m~G��8��2E0�Ń�^sƽ�Fx��-tƳn�Ɏ��IN�iln��a�uO�B�1��/�7$�&�E��6�=E���J!�h
�C**yEh5�)�v���b�dgPO�&K�SՑ�������8� k��+�W�(�/	�H}���=+�c���\t�.�#cw��FnAy���e�@��QV���n�%k�+YNNN�LB�G`���������T��8��2u��X�٘ %ZJ�9>@������T]�q�O�!ն��\I��׿�!f�u��:zz���|����z{��[�.�����g�;9��)���1k��g&ݹ����J/�h2�i-���*��߲:&�<��$E�`>��3䃽�͞�3�0��S�\�d���;�� �e�s�������s�V��}������Z�)��*t�����p6h��WR�ۆi*�*��;Ե7��nt�2�-�R-1"_�ߖ�2�K�U��ɓ�B�[oI���`��_�ހ��!�����G��N9I>��C�u��{�����ug��^�v�3C�s�#6f�ӓ��ˍ�Ãr&c����SP�Oٞl�q�j�g4���4�����C�����Ԍ���Wd�-Fl츠�}�����W�ׁ��G���s����y���4֪���D=E��ZFK����G ��z�-�ʾ:UI��qq�9���ޓ?�Mg�N�)J�<��)��9��2��æ{_��o�戶��[#$_�2'ҁ���>7Fmw�F>�{�WSe���[�#�Q��eہ�Ğ'@]����ƭ�[Ϯ�U������S#����t���'���	<A� ���KT���.O�vAɮ�eɎhA� ��`�孞������O�͂��_��\��4I�m\������N����Zk+��-���\�@e��w�m��S�≱���bD�y��ZiF�{�U>�g=���>��dm�o
ߎT��(Η9J�����Ǵ�����읍~hq?н�Ys%�uSi/���;�_�ja�$´��"$��L���s�
/VR�x���&X|샰����u;(=�J�<&��8]I�fʞ񩆛dʙq�x�*dcr�]c!��"e���w�y��r�,�[�*��~'�	r�zG���&?���?a���~�_YsN#����N	X^�7�Ջ�B]r�F�iQ �����,`�qḌL�c|?�s���ժb
��=�l�X�}��*��*�EQY���	>���x:N'��+��C�~���꿍C���#-���B�*�m-aĉ�U�]Q,�A��+y��:_K����,aC�	`^��:���'p �`��������.�b���y<GW�h�/B~|"�[�+J��{�k��Xq��*��&>�rգ+�}��af�0�J;ӡ3��W�$��P�)��0��%�d�vJ���M<��5��%پw�Tdڛ�Ax1����OQ0�K�#�G�[�5��ȇ���p�����6�������B˦VBb��m��.|`8ޘ�R���w��*W��B��#���ds^��!���|@zrZ�;��L5���zpn��$�Y9qs��[��(&��Y�Ya�\��om"ÿ�C���L����A���"�p�1r}��H�q�!w��("�C�D�A��b�w�� �ng�[����ݠ�4
����d)�#�^C��m����V}\O�]�� F��%:0�)��p65vB1�(]�\�H�(�\j0dקCbLw��]��u:=+�.j�P<d֬�,�-F�=~.2V�h��S�����a�'�]Y�(���NuA��~�Uջ��Vo�cr1:��eɩO>?�㹀\M�S["�+�� ˹.��$��C`�9��#x4şk��RQ'A�*]�Y�s������9����uҷ,�<���y.� �V�P�H�����\�����i�˜Ύ?�����w����Խ���}o�A�Ӓ��y�����(�~��]+!V�����풣Ϻ'�0�}�\yF��!l[=��5.�{$K��z�;����	O�y���R=<�)���yo���6?x�J�3�y�Q�\RBψH�Z/ۼ9���o�I^�qM(�'�_T�����i��#� !�@?𤺶���G�k)�ٛ��I6Lrz������p�Ʉ���U�-;ldĴ+Hq�,�r�0py��Pd3�遾��Ϟ}`�i�o����g�8�N��"�w�@N�߯\[�Ϧ��X=t0��oot��X !��GA�P�Y*��Y"v�������*��x嶫���-��廮;��H ��%g�c��%�y���6d��� @�}��>L��������������7��ïn����ѫ��WR���	_2���:��޹��o_���/��;LWI�XI��]|�@s�νv�n��%�/�E�{��3
���uA�S�#�I�����M�u٫�\���d��x��M���y� ƶ߾�¯s,��8�N@������x�$H]y��z����鞤Qq��q�^=�so�nq�/W߿�k�t��8{�<N�y�_;���W�w��r���<��o�Vi�oũw��Ի�p��8�>���0��e���S�y�v_=�t��q���aƟx�,�_������c8��Ey�<�:��7N`�kG�c�m�yD�-o�_o���wNa�����a4�v�71|�o���7���#��
A��~�9��K��51]�iy����[�p��I�0���a4�ކ���A���MU��T_ߏʫ-(��W���>T_cܕf��o@��d�P�9Q�ܓU���F��Z��S*>_�ҋ���6��%mH\��f�]jRe�Oՠ���k@��:�>R���U�8��i�(&�f�T ����v���~T5�"�2)u��u�;�bבr�:T��i���'��)�(�Gl�v$��Ď�5ӷ� B�NϢ`儣|?x6=�ɝ�Ay@}�B�/ Jׇ�U@�8�%YQqB�by���HD�,����Jc?����L#��q#�\C	���n;�v zO"B˷(�� �V�.	�U[UC�OB�2�?��-_�������̼��W��0B�H�4�*q2�J��۩�ц$6���|���ψ�8�Z	�A���`�.}kB�G u |�IwĺLgl�u�Gy �[�{cP	�Rlʑyå�O��ȭ$��"��B� ��̄V���*ޕ��pxd�7;�	/.qn�2��_�z��C{c���6b�N�i�:�՟�ٳgb��`��l�ΰ ,�b��,�#�͙����3�=f,�3=�� ���f[�* �'l�ؤf��"��R�)~P[��ʵ2����5̍m0}�A�������a�d����j1���̱]��������Bذ-C#K���Ș�J�L�#���YB�#/� ���4~,z�n��� �
���ٍ�C�ٟ��n�=��p�=����ڙx<�q��m�s���㾩��KdF���w;	�m���ME��V`T33�ɌiG���o�t�F�mKp#+��ނ��ߴ@8���c�����l�J�+��ƋIԎ��w t�t�B�΍XC��HW �y����A\z�W����	��ݿ��y�L{��'@EP���FZi��E6����&I���_���4�D׾��/ �$�n��~�!I����2�ն��¿�>�]�C���K��^jo8��ۯ4>���^�;���c\�d�@��FJ��y[�Ǵ�)�̦�n ������?�R#�� @��%�WY�Ա�n3^�T>	�2��8����7��{�?|Ex�-ˎ���4� e��;m�7���H�߾�������w?}��ŗ�X���h���Ʋ�H|�i��GJ^� �������KɟА��>��C���{�>���>i�ж�K���r�o�������@��7��ӯ?V�~��94˚d?��;���������/��W���/>Ʒ_D���1,����3]�x}�����q_~�!���f�E�H>������a������=��Y���oY�/j\��<���2ޒG��;����*��g4�[����/�J=�<b]r�%ߧ������}�.������=|�q�����w�Ґ�X��/?��L���I#��f�/���� e���?S�M��>��`���k�+���S������{����歛������oJh��K��mB��o��#��c���g���/�7��[12sC��9��ωo?T��������-����p���4ޯ*��͋wt�K4�i�����M���U�շ�(����ִ7?~�.�Hfz��go�n}�����dܛ�����o@�:���>ᾲ>����EB��z�4μzg��o^[,G]{�:nHn����Pᛟ�쇯�һWp��t^D:��>����å�Yﻧq�Ӹ��E�����kJ�~F�����M\��.z?�X}tI�<�C��8G9+ ��)���K��Chy���?��1� <��Eh{��Dx9��)B�QB�B�1}���N "��|�Nb�=��9�u�u����Q�g�Co��$�ґ�O���W�(�}��q���s�u������gp�ud_:�=�v��Gh�{��q��	J���~�K? ��Rn���� �(Q���Q�ԉ�.�����wܓ��T_�2���7՟7N*������Q�ӌ��{�eNs��}rU�)�Rf�k��GP� �r���f�U�x���{FI��x�[r�T���h���������uU�R�|� *p�7���}(|���"�Jr.�#�R2/�"�|�R�=ȺXG�+��ۃ��_�t���J��O�"�l�E�+mU�
��.Bȩ"冞)F��B��+B��<x̈́��tx�T~�Cip?��t=���8�#J�'rnIVr;����|1�1	���e�Nx�����u ��ӽ����-��:��#Y�>�	���g��ri��Ɲp ��7n,�q@�a��2��:���1=��T>��'y��qj"P4��vEnͻ�ژ	��8եa�]�\���t�lGA��߾��G���^ApA2^��g�C�\Q4^&P��Nd�$��&��z;<��Y���8�0~Gsv�MCTi,�r�����|Q�@]s��F�t���'���=	�"�<���KfP	���O�F��i`4�$~y!pM��.O�"�Y�� B���D`��@�[�M�T$!S��3��W�@�4e�5�2�<����2ތ�`}lۋe$,n��W��0�'�JD˅h�j�-�;�ʲ]#i7�~+�kc��Q�T8�3^�
ByU |�9�7�
�d�3�A������1�^��<o���OC��|��@B]�.�%2�f��B�y���M���zz�G��0b�P> �L���1,��u6��3֖f�23Q����l��ޞ j�G-���N8o'7L9N-�]<{�Z��?�m�ӵ���L���v��9�1����5�S7���V0ѵ���%t�"�f`���t����F�2р0jS�5ҟ��S�ԩF00����L(�:��F�����`��YX�qV;9�l����C�ǐj9n7�C����v\y9Q���ї.�h��pX=b����`޺�X�O�=��.p�q��L	�
|n eX�����<��Ѝ�wCf��̨̈���d	�<�&m����OD�GH�5�+;��;��>x"�E<����Z�����\K�\��)�,��@7m_��%���
���~�m�ӄi<+i���[�Y��h/�Z�$|����u�w�#���e��R����A��8����ϒ����u}���ְ�?
�@�\ɗ4x?��C�O��cԟ�x������}K`��#|��G��>>��|�#���_⫟>�����}ͺ�U��?��~�J��_��1N�F�G4p���?4�&�U|��~�
���|?� ����������q닷��'4Xi����7��/���_�{�/�E�V�U��OR�p��i\|���wW޽����0�q
���;4�o]���i2�����p7>��Wh_~�*w����1�?��7>o~�^��,aiC�^d}WŠf����$�IqϿyg^�˼ט�,�z���[�p�U�L��]���oM��اWU�$���7p��s8��\��*�|z�>��3�Ш}����νw��[z�;r���5z����d�O5��L����KqRf%���Q�o� �Nc��-�+�q��8�3o���[��w9n����Wq�=��]���4�>�Bi�N�o��l�������i�t ����F��E�T�A��ZT3\s�-Wb���J-����>Ԝ�G��:ԝeٳ{�x���ᄴ���.����p�}8���w/���}tUş��:N�wGߖك��{�0�D3�}2� 3���~��qM���
�zy?�$��i�.e�\hF�E��W���J��3/��f1�i�6�Xo|�8u-4�[�`�A|��9��K���7h���}����4��Ѩ�Oc[�G	!Gi�K����-����x����I���&�%}��H�QB��/���g�p����>���B�咫M(�܀�+M(��寴P�PAռ~5�Qtk	EuܗZ���%\Oc���y�{��� �N�Pz��}p?��C�\�A�� ����L?��������D�~!��i�4���0���퓪n�������!u�D�U��aT�y{�9�Z�_����Գ�&i�Kh��*�=�ҷ�荃J%oB٭�(��ܥ�����Ux�����#(� ��jA��M(|�0
ߥ���:��� �}�~����E��&��ڈ�7��r9⯔#�j%�]�B�+5�~�Ji��j$ߨEʫ�:�|�;n�#�z�2}�J��^�P��?�j5���re�.U#�B".T"�b���I8�L)�O� �\�
��-C�I����S�*O8���W(����z�!���W� �J"/�^�-q�Lf}��s����c����8��#/� �e�X>�z=b��h�I;ү�E�_їjT|��=�r���D{����"�&�*Sn$ێ� �-Sq"����?Q� �[ �)�t1"e\�P�O�¾�)A��2�����bx�.�ǉ|x�*�'�~<.G��D �L�ZM�z�)Ii�l�l=Akl��u�����4���j�x�V<R�e4�.���(,)��b��%4���g��x�f��Sz�,�mZ\����-�]��(�*��̲p�VD���"I�S�9u�[��p��ƹȬ8 F�>0��q�/L
�Tz�<�e!�,�){ɧ���T��x���E��rMs}`Nв,
�UI0�)q�	X��+b\q��ę���l�J��Y.��?�0���%��8B�I�/��ܡ���d�(W꒴i�\���
�L/�f���oXg��67��ܟ?'�B/l-L�V!jަE�)-�Oi%���-l��1� ��u��u=��8�(͕e=07�����ڜ �!�EAWf��Jb��M��%��%��W�kP�6 ����xI�ȕy\��V��E��*�'�S���� &��;>��p��K�<s	V�
�|�'�V �3�� ��eD]"�j��[�l��}�6�	�Ҏ�׃�����֋e]�.�`w�����{�|���?B�U�X� h04�<��[Q�HH�N�m��:E��8�#`W
|��|�<+�]�|���ff�D]���ֻ�y�96eA,BpW�_J���J�o�eC�<w=K9���sEn���T�j�7V������= ���ǰq򲡁>v(F����&��� v��0w�=f�Y��Pz�`en�%�����exd�|,�9/X�Ȁ`||�=l	���q���v��]�y6�4 :s>at��Ok¦��\Z��,��w`T�f4H�u�1m��Pc� �,�o��}�M�4W�)Pj�tc�;� ��g�V�01��ߤu�B=:u��jM������ᅗ0�0=Hk,z�� T��>ػ����=ѳgO�����=�~�{b���_i�E�b�F{,�zk	l�%O��PyQT����B��� ��am��r%N�vhg �>5 J@�w@צ;`u��7��ذ��̍�7T��.���"h%��\�bW���xy�Z�3�Pϕ�6�u�@7$�Uo��g@���q�"􇟾Ǘ_�O>�J0��c��ћ�����+8�荳��38M�y�4u�����5��.A�y_��u�W�'4|����M���-�����a��O�	��/�����>�}�1>�8�?���;�����w?���|���a���>��ƿ���x��w�������*M�H�[܏W߹��ߗ%T�����Ｂ�)���;��ç��P���4ٯ��Fh�J��N�y�߽N����%�����p��9��q�	=�o����9Vo�#dpܨ�o2��Pt�u�r�ԑ��r��K�p��p���*�a�<��<���Wp�0r��L�B���e����RK�$|�#�҇�q�v�U���8��S�,�h�;gU��ۧ���7�����P����yͅ&�M����7���AT�ҟKM(�؈�(=_�ѹ:�\ۧ�I\1�U�ﹾ�,#�������jo��W(�5��#��2UW�5e�r��ʭ�"jVu�x�EҪ���rR_[?��)y��*���)��%7�Q�
��ܯ�Y窑}�y��sa2�T"�t��#�R-r/֢�
��UB�넦�пO��6 �\�ʟ~F#)�q�i�ʑz��O���̳U�[����c��W�����(}�w�o�l7�B5��U"��<�/���嚐}��r���'��c���Wj�u�����8q%�M�'��E�4���l����I4D�ϖ �\��o�H���14Hō=Y�x�	gKUZ�_�'Ӹ���g�U�h�Jz�Bl9Y�h�Q�r�?�4����P�8�D����̥�}�QTȉ�B8�l؉��l0��?�yG~��K��@��,���e�<��Q�v�.�+m�����-��	!	���a�PQg�T]ҏ�Ӭ�L�r��e������dx��<�^�Ri�g#�$�*�?��?���!g�	.�>��|yLc�~�X�D�h�N�xJ�������9>	*�_[Y�ϑ�рwmNf�v1��fM|�f�z%�� ��ԭ�s�ݏg)y��#@d����u:>g����xp�ܙ�r2����v�q���y>�������r<�Gֵ�h�MG���vR;��E`$/4����mxq�v��V�O�-��\S�m��34�������>�k��0����X<ִ��Wz�%+�oÊ����D<��%-qX������`"��ۊ�{c0�!�u�ʝ[��0�e[��[�hnS<f���~��ر�Y{b�'���x�oN�?vw�'�2�.�v],�$?��3�����(�l�mM4lY���7�i����h�-؛��-�0�is�ώuK�f�V��FꬉR}�<��\K<��e��'�U�J6�a�θ̪��%�kF��+�cYA7R�I؆mH�����˦>��k��ŵ�q����\��0�7DÄm�M�1�4���y}���eٸMq0��s��w�>�ϐc+��Q\I3���2ۻ�<�D�<�뷪4C�z{�@�2f��`�s˘ch�6x�9����ԧخ!�'�C;`|p;�'B�c7�)�.鰿����"����h�&��t�O�M�=��t��TB�NMt����i�����јV�4�c�_˶�J��H�aI��k�i<^S+hȷS[�.[�Pe�V�C� 2�,Lŷ��ư�܄�nP
=��ք j���Ÿ��Wx��!~��[ױ.��z��	����%��/#��º0 �+��DYV|W0���V�}�~C�,?B#!I ��u��.�ߙu%<;�� ub�K�B�	�2#�N(�߫�&\*�����e�<�r%��_f5>��|�A� y�nuB�l��	�1p�e�lû$�"\�-�<�lˉm�2��Ȱ�"W��aԙuK�Wy4�0�2[K�ުfN}J�Բ݀�-�9�� p|F����+ �-Kd�8��� ZEЬ�K�6�x( ݘ���PD�ۆ~N�gV���C`	�ۑ��E?߁�u��/ԫ� *yY�,��,��w�]�ūa����u��?�Gbĸ!?y,��-�	0�1�݂�X�l!�/��Y30s��_��=�V�]6w.��[H���%��ղ[+#���Y�-lLl`kf�E���x�R,��Lg.���B�|��3���r.A�^#��f.���BX�ȋ�fb�>��)��:�0Ե��̠H��>e�	���3M���b"S3¬�XY�������>�5��xz�j̴��0p�h�:��8	����F���^=г_7�� �N����������B�x:�9T�����X,�n��
|��>��:a}�,�u�+ ��\Y��J)�Y�lgl�q�̀@�SS���1�w@����K�\R|[�e�+�j�����m]�����M�ש�����0��rz��k8|�j5�����I4�<AC��4����S���i4�~�:��7O���3hz�8�E��#�m�q�,����8��9�)K���(!��UBץ��#8|���¼��\:H�0�� t��r��g����>�|�Waߵ����1���&[�h��M,�x� w��`}׏)IX�$���Sha�jY�I��%K��a?����W����~��o	�ߠ��	�s_�^;��׏��aqU����7O�� W��)��:��7����({� �	D���O�0\��>BL�;<WQt�I�@M�'�l5�9EL+��e�t�����2o1�H�B�Q`t���J#��7 �@�J`� x�2v]�F��^�A��J$�-G��R�d��+{�̴�K�*��bUk�I̛x�ۮ$.�O�\�q�(C�Ä�0ǡ�	T��#4���!�����K�4�	b<����Lx�D��K�i����ߍ@����U�k�v��W�.�e(�:��:;��T�!��єϽ�:�� �a�h��a�YJRV�%��"��	BQ�y�!��+�L�s��p=�.���(!�X&|i��+�q/��w���M�\����I�ȃy\��M��Tr���G3�&K�dI�D��ܒ'B�]:��54��r6I��y�S�J.'		'	�!w��;�ȉp��h:6��S�f�4�_O0�, ��l$����+i�t`'^�Q�4��h�=B���<wp�=��Gh$=A��i�����ѷ�*Ki����GY�)��C;��H
�ݿ]��Dc�Moې�
w�i�>��Ghl>JcK�'Z���<t�
/�q&y�X�W����MѮ4�i�.b���x�/�!�0�	��a��Y�Q��R���6R��Ѐ|��[��]̺�s?e?���	���-��aAfI�,&�,%�<| �h&�H�⦘;Z���do,�[��1꣔�у��;�đx�0���6ֱ�u$`1ۙOCu�î2�t6la�hƅ��<�4�ӈ]�>.�A���g��4`2m)��4�%n��ߞ�=]���1��m�^BJc4�q?f�6��	"�g�	#lR��0κ!�̈́����,�v-[T��ڢ d���3C��K�Xf�ඡf�39f�O�L�ef�V�"0��&ʚPЦO�C�`��9���)��kq��q��p���	�#[1�l2,���I�K���8%t�Q� s4��Y^�P"&s?tx���PR�ǒ0���{�`B��q�S��<F'�a|2Y���w���.��O��	����09�~P�p�$�ى�ψ燤KXdzLʳ�#Iܟ�mmJ��'v���m�_���2M���7z��Q����~h+�-���$�{8:<�uن�"��>KXd�}29���u8>Sy���=�-�g[���A{_���O�X�މlC���H�'٧S;1�H&�8I�$�/yƳ���۠�Qܗ	��9�ٗ��R1�c5�@��D����S���IG5��/Sym�9�]^c�O���t�΀!]�c����yv(M��>��)�O��b?�������R�V�V���|�a����D��RF��sU���;a��s|?�ڔ�A�x]�(u�3:��c�R��˴q�6����5��D��nL����D��������Iq�x�G`����-�f�8^�G>G<�6G�Z>��ӱ�7�&
c�#1����L�Fw
?��0�x����aQ��nƦ�t���s|���,���Æ�D�F8�$��e!�*���R?h���EU1XQ�����B&fZ���4�8�9�L_x����̧f�ϝ��#�I %�I��D:3�A҅��@8u"��]��5G`U��.5���8׼ 8���1ӇK��gOU[˂P�F#X��,#��"�pF��'�½H^�7����%P\����X�z�S�	ě�7G�əe6�%�ʼ��O UfH�	�����)�"�F*ɳ���p�}���}4����G�yM�*g�
@}�^��� ��!��{�O��\O8�x��R	�6���V���LV�z��OF�tlmJD8!4�� �},��R�Q��0��ވy/χ�2s��5���&�����C�l:&Nӂ���z�i,xt1?��=�8�|�)<�ܓx���X�t�.^�G�-Q ��R�Ѕx|�̈.�R��Xh;� *υ
�Zc��L�-$�.�cK�����picn�dM@�!�p���dlg��|���+7��/as�$��2�0ҷ&��ӵ���L2lHwƌ�X��	̚�zz�04�R :m�fX�b�Ű����:�<� �[O/<��s�jn��Ӧ�ߨ��6������z �z?�����G<��Sa�%n���c��28fy�������T�~"ǡ��
��<]�� �.��
\�2M�B���@�,Ͻ[�r�M���l���p���qOŖ=;\����It��/8'@��Ux>f^�J��F�LZ��/�\�B��>�����n��vnFtkz�]?�?� ��/Dҡ|���x������J=�_�C��Z�]�B �����R���U�b.1��K�JDZ��W �\���_�öM�F8�?[����T�����J��=S��K�j��6�G �#��1>�l1b�a�-��o�%��J(�V��k{�9��+�\	(ۯT����e�r��R!(V��Ks�qg�q� ��(�h�Ƹ��ԙB�m�}O���X�r%ޟy��K��<W �Ep��/F��b�+��`
ֵ������_���e		��`þdl��~o�6n��u�xqO������e��>ֵ���<s`�&$<}p�F��>A����4f���'F�R��h�>̼����`��K-a^q񂴀��|��i�/�Q��7����M��Y�7�sy����і��,��x��o��h<����ڞ��=o��h�,��0g_�h�ΦA'�Y��PXׅ+�mS4�b0���<������}-d�粟�	��ib���L�R�vo���g�o�����E����3���	��؅��O$�q�5q������q��q��}��1Xr�0t*KF86ү6-lu�b�h��ڎ94@f���<.�i���Zt,�%S)Xȋ�<�f�fb�7�~�'��q]|������@,8�֬Ӭ9Ƅ����՜c�1��(vGv���(3y����쏧a���=���<���|�wp�N�=�O�C3����S1�d*L�w=`z�۔�a.��x̘ϔ��`�9���7�8�t��?���>��J���ݘ�6̎$Ü�j�z-e_�Kz�����\��7�7cS�K�Ђ�剴�*�әJ�4(���zU4:�=iG�%}��w�ī4�I^+���\&L��K0>�C�z
��&�2���B�/fÜ��M��O�S'u��K����o~���2��t�p,N�!��l��k�<F���K�>!�3�a��:M�M�>�M���z�����K��.L?�
j��L�&�"�M>Ic�x��d��4��ʺ����a�%�3�I�/�R�gvQ���~Lᾊį��[�Q�N�R� �S��I���I�[���4��n��ɱM�j�&s�E�DH��1�H��pgRy�i"�W�cߙ��8��5�e���	o�	��R�D���&0n��mw��x�� uH{'v0�`F��q�z!��QcXv4�h�1����A����ҿqڱG��Ac/��I_�)��$�ƕ�������&��I<���X��X��޻��I�*y�����I�k$m������^��K>^�%�8���hJ`u,�c	����J�e�����1j���p�s�y�C�k���F����M�@���e_jb1yO���:���t��<�1�W�;��)YI(��¦5�i�k#0�&ë�0��9�"�˃1� �U
-��8j�	PSc�Żp��O�ͯ��H\��c��N���a��Z�@G{c|��}1�0�h~(������>p�CX��1�U	(�T��@�#(�C� ��p��@����9+k	�����Fʁ��A8����aO�h��Gܘ�A��M8vc{�lϷ(����ry�m�*v!�b'�+��[��P�n6�	fN�!���ea�j�!�k3e։ ZH �ǆ\?%I�8�"�v�̈����*�ԗp�SOB��I�wy$����_� �Y�!�=�������e>p+��G��k�	�A�#����|,C����}�ȹX��=	�mډ��m�m؆�©�ب\`��>Px!�}��/��0t���b��Q��a5�s���v�L��2���b��z<J贴�I%`�x�?��?��Y�9s����
6�l[[<��<�h9��ÂY���#��Z��k�g��;B�<,[�(�X��g��٘IYY,����&ƄcjΜ�X��	,^�6�U{��Z��hLM�ai��Z c#�����fНn���V`��00����e���`*oܝ�&f6��c�	S�ahn�E�<���7a銧0���ƏA���Р���>=�`��x�oO<��AB��;�;��Fc�c�X���ݼ�Ƴ[���8>�2[N�/�U/���r]_��sM�3V8au�3�T��nɳ��eCwɃ��\�)���6Í�D�ޝ�ޓ��(8��bs��z�s�?��X�g�����Ux6����� �+	�/�"|�Z��)k�� ��@�j��L�\E�C�f8�t@�;�����ӑs��ݐ�`~��7&a%�i%�����y��I�34`�����F��	�Χh<?M��)�OR+h�?ּ�4��Q�O1�Y)O�w�R���$��'i�����x�}�H�E�	�)�=IXXAc�qԒ�I���`y�x
���.�+2�x�~X���^��!�4���i�>CXXqx%8H��L�|"iW�K�#�i,�x/��_q���>���`.o
�P�~��fSs��P`�B�ٿUɎ`5Gf"x���<�$%�fof2m�!���%��@<�9�Ǟ���a�ŬFY��\�(;joB��f�zLk�`ȋ�au0�kB`Z�,�x!��>��f7�7,k�"�Y��%��Bĸ6��N3�IC���hgɲ��7f�Qc��ǰ>R�F�Fu���29� ݖhLo����X��߂i�Og������/��`t(�y�(���V�c�?�*Ǻ�av,���H�I��Ŕ�1%Ȋߊ��,�6<d�C�rh(�s|9�F��Ä��xX�,y�
T�i�g��t�d��;B�A���v��NPaYB���3c�t-y<�����eY�8�K�#6���6�Qb��,i�Y����9-�%�ڰ2�3���,��V�싄m	�F,�w��G��<��Ǳ�RFlׄ�`�sΔ}W�+$4��d��j�r�$M�`i���L©?�39�6���$d��,	=F4ئ�]~>��(��}�aD`0�X�����4��o�}2�a�Q�4^�i��@7��OY�F����1��nH	LY\�&�e�|*�sTaɈ�Ș������x	�ŵ�(	K��iKo��i6��8ϸ{Ȑ d�2"���I��2���<�5`�6��t%l��,/aS��ԣI��������"A��2��>��G��#��Φvt;H��L�(=�����1M�;5]�p{M���%H	��x
|jS�:�Y�����<�?���AStu�i<��#��$� �3�l�D�群 �����e:j"��Q��;�*�zd<d\T���a��^Pw����ؓ;�@��?֯i��F��6 'y�j�S}l��*��V��(�Q���hJ�����%�Jx,���1��Q�[�F���^ *���j6U���n?�$���҇1���~,�=�Z� �/���
T��=z,�cx�������,��c�h��L�h�kGцݤL�����&�j��$jb=�ȱ�KVG�ΑtE�����6�x�6�iӌ�z	$�b�E�C�f�I�,�E�[�	k���Owb�F2�9�p9��9��� B瀲 *C�0��Ȋ i�1<>�c6amq2.|�)>�o�W�]��}8�쀮��zaj��@	�c�ܡ��	[B���6 u*G����ڐBcx;�~jf��LXsf�� T�S\� 8>3�9+ <	��<���( ��GN0|YΏ��!���K�d;
x��U� �A~"%�"QU�_����\$֧"f�Nx�`gy��`l 0Y^ ӵ$�Y�,/�����LO�%�n"�n0�~�g{�V�r��0���*�GI8��wy�E( ��茀?����$
ԧ&X=��Q�Ϻ|��*>���>7<<y�dӫ4D��(v��:��-M;�K�b��Q{�bKm,�/�<��%~� �:\�+4���l�j�-5��3,~n!<6��[��r:�f����ֆ0�2��-����6�9�s��\j��x����e?6f��`�<{,[��̇��,̳����1�n.,MX��7��im6���K���cau��\�X�?�~�
���Ԉ :{AӖp:O>�
�=�"���`���#/a��ga5c������0з���<���xLL�g���N�j�ً��ܿ�00�¸I�0E�/o،��h�/_�1Ӧ��葄���/��{�[�^�֧� z� C��x��lX��.�1�m)�>�<?��Z�Q gB�#?;�2�Bha; ��� �y8�35��덭-�� �[�;���	�$Y��"7>W�٨�x~�:��x� ��~�'Df!)7�O��O��ErSB�dbө,<w!�����XF-=���4���YB�f݅�|�h�̣�"�K����9��۟H��g�".q��6oR�9�4�7'KB��1�Ƿ���1}4���v̢��H�u��=�7�h�y���M��P<f��4�-�,�DVGU��Yڪd�vlئ�mj�����8�7M�m�?��`|�0�6P0��M����Q Aɘ�`r��r2���NXP�w�0�SƙP�2ސqF4D�4
LX���d�����\���W��i@I>�o�m
n��X��Lx�T�T\�Ð}�g_e��tj�,�b���O"Y5�7q=��t��4�ѥ_�F�ۖ������	�su��ܷ	<~�٧	��4j]f5��Ж�9�S�,��7��9����)ܧ�L�8��4���I:�,�.Y�e��A��H��,p4�F�x�He�RSi|����te&�P�Ki���Ԁ�}�Ʊ���t���g��ǾLU}d�(��O�ǻ%q:<��r�p_d�&��1,�>����ҧ�#K���m[�gJ�Z$a��6ϯ�<����Of�I<�&SSy����)]��t���#���4m{J�HX���GcX���4��[%}�16��͐�s}�w�X�6���;�}w
��)�<N����w��~�1��xGi�30��0�T�>�z(�9�a�t6ʥ�.Dm�j�7�}S�)���u�ֲ�DJ���w:!M�{>��<�$�w�$�yڅt��:�nq�H/fB_f�f(�� U3;)j�TI��� ����� 3�
圐���S�BgZ�$��fVR�ֱ�[��ʎ��u|�p�'��v&m^��Yw�&�J��0�m)�θ	�Of� 	41ܙh����U	�q��/u�ۙ��̵I��3i	dݏ���z;�R�� ��/�EI����tWۭ����gt���tT��5M��̭���ҕ�8^?����^2�8��E�rۓvǱ� �޳��r��#|�i�iu�]�GJP���H�#y��Q�̦�m틚�m����sE�ؐY�1�OB�8^�G��ötJ���}r�j�Հ%��
&	�2�)3�#��`X��� �� '��2�)���	�c�D�ΑP�(��i��Vj:��	�u ��J5[�� %@ڿ�40����hL`Y-�Ϻ$~Asl}$ۈ�����+3��Jx|M$�L>�f<E�����L�$�V�ߕQ^�!���0 ����TcP�?��)����c,k|4΢$���S|J���@����)����b?�)�fw�fy�.' �ޞ��Q �\���$�5$#�:�Qp�	TKc�D�re���B�J�t�
��t?����w�L?8��]��f�����=��HX�L�����3�L+���AXE��Sf��l9��U �X>Rg#�,N2���u܏��ʍ���YfD�dyc��tw��F�]��|�u"��:���9��]�I-�~��J��!J Ո�YM�	W ��2�Y�1*��k�'��(���	�^�cy��{Q ��\��=q��Px�!�!��x�G!��Q<gK�S� Խ�u�;�ݸ���a���=����L;S�[��tt����Tf�057���̭Ma9��sg�~�fϷ��G��ٕO㹗���O?�e�.��l¨�fͲ���l̝CX�;��3ag56�3`mj��tţOROa��eX4o�ҲE��e�a!��������=-,����Ob�g`g�0�
�s���%07[H�}K?O`}��am��к� jO�as`e=ړ�1o�2<��s���=SB�X��Z�
���xy�&�,����'����/%����,}{�{��P�?�gA�L���9���#��v.�z���&��C��˟x7˛o��C
B]���k�*��?�����eT��ؐስ��F�&"�2À��j TfA@�'��~	�@_�J�L�� uIތ�����ç���g���7��2��|6���y�j��,��x��l.f��F�hƅ4%Kbm�Ȝ���"�]ʸ+�H�����.q	a�>O�0w��v�pKV��q�EY��M�c�Ԍ��,<�
�ӻ[�
C�mĺX�>t	�+��KC�-N�kț�'c��	��.e����?�B �qNH�g>�*Z�K�]��y�Ӏ�~}�.�Ez�{:o�J�W@C$a=�7��[[�n���Ӹ����y�a�SY��	M��x*o�:lk���thL�а�¶�0<��&SڼOb�	�D�w"۝�}O(��K�c\��2��O\���i�x�Q���F�c��;��b{bh�q)a�.���~�z��J�����k�Ư��D��'&%�M�`
�q'�eM��I#�'�&�Md�	�G$���$�M#���7�m�F�?�8Vc�W�|��EM�qa�ĝ$mR�ih�g]���1�b~���|��<'d��4��9NƊ�YG��ưָ̘Q�q��%^��~H��$L��0�I42%N�z	��a3J�����sF�fh���5���|�2�b��~j�{�m�c�d�	�gx��'����%�,�1����M⾋+�Sؖh25^�x�E���kI�%p�f���N�ǳ���xRN�ϔ��8jq<'���T�����d^?ĕ��4m^#���D������}D$eT���I�Ʉ!�W#�k��� �3��&U��j��	�I�&s$,��fi��l���!AQ���%N���k��3{)�)�/�ɰ���#j���:E
|�G��c����>��N`���Z��s�~$���I��'��N%�j�yLT�?�r����w2�k*�&3rcx�ư���l]�Ƌ��C
�8�Rf�"���ߣ1�N���z�xN�����婱�׶>ݑı=�*�ϭ T�����irm����pd'��s{���L�v";���_�I�������Fu�����.VG�LG	h
T�lMN�~ �:���uI�ow ��Î�/#B'�:j�G���{hľػ4�%ed),5�M�������!{	����4�6G.G$G��/�Iw$RS�u�.5*����
@et��j.%},�N \NdYm�5��SXF[��0��I�s|]FFFJ>E��_A���j�&���q�ֽ�7S��0�b�݊(����Њ$��!���
��� §?�h TfD��Ƅ�0�ߦ �3�����/>�WiLB7B� �M#wL�'�e�bx�fLIuƬL_<J�[��2|�J�� ����DDe<�	�򌧓�\��w*��c&A0�Wi3%Kk;J�딗�|��?!
L7f�)?� �zP	��^�;�2�'��݃���e����o�!�t"jb����3h��,jA �g�F�4�٪�inJ�_�� T�S�/�r��Ol�.�X�*���J�s)&�F�KC�UB��@h��ϮxT�2\o��(�R/��xyW!pO�Z�)/�+�,�,����hI��T���m�DC�ǲ��OO�~l3��Ū�����LX=l����Ƽe��3ג�hccL�>�t'��Df�0�ׁ��t�f�6f�����B;���Ǌ����/bզUxn�K��t1̬,�o$ k��b��,M�1�fH^�/~+Y�'�?�'F�����*<��������%̍���a5c!��a�����K�X��9��"Lי=��0ЛC��z��=�����1cll��\���1l�i�9���h񣰲����l��B̘EP�i���z�����l[����#�6�ǀ>P�ڷ;�@���0��c��2,�|vN�xس��4�NfA��O($XnV/#r��"W�2�9lv&��wf@��̀�V�"�4>9�ͷۙ'�N;}�l�Z<��<��\����. ]�c=6o� ��n�L�̀��;���D&����yW21�R6l(k��b,�R/y�(ft��f�w9&�e��,K�#E�6���;aYn7�f�tx�	4M���piL�4<�2GR0�x:,����X�)�c�aư�	�w��g��v��X
���R2�G^��Ǜ�o���I�1��ZJ�ƾ�vC�kD�Ř7{qM�Of%lКG�0됗,����%��ۊ���N�d��!�ed=G�X��6��}�U~��Db^�Mߟ ]�,a���:R�Q8������cpXړe����C,O�Ȁy���i�oZk���6��ze���`��lIq�ߨ����o��F�1�͐hKk36D#Ĉ��2J�7�V}���46یI-����� 4��#@�g��lҝľ�33"m��� B� �\�f��'a�_#�7�c.��Ld�,�|�0 �l'R�)�t����a�pB��֨����_���5���qԒ�y���?��Q�c<��|ۑ�q��Xۑ�i���P��Ibx�F#�MnKI3�L�/F��i��'iw�g"�Cܶ>(1M�2�)Ǖq�9��Z�ǲ��9^�y^L�y3�牼tC�CM � � L�h�Q��H ��#p�%�!�&�n-#_ �g�{�I�)�	3�嫙��<���ra� 0Ϗ�<dvT�]������w+�-�[iO�$] w:�E�r&�*U-�Y=�m�v�h���9.�(闪�]��x�J�i"�I�:�i�r��$ &c+�H��z.U�6N��C3+��֙J�li*�v�t�S����*i'a�MIX�Z��_^O��nR�˔V��H��:�s�P8�?�<�r|�ɱ� ����:Ɵ�9�z�1�X�z����Q���ֺ&��D�����v[��i!T������,���4�������Ԭ�=��k[f��NG�]��K�m���?������ڮ�m�^�>˵��:-����۫���^y���(yq?�����r}(x������T[��8iS�k�m׶���;��{h�A��a�N�z�Jx�������6��"�ScHu��VV��s�� ��V�$pv�0����L��R S T\���O�X�2�@'���Bfu8F��KY
+3��#�4�)ee���ʬ�<��%����O5p	�
TP	�����3��i����8�6�aau�̜�s���	�7�m#���+}�&4L)��d����tx-�Wf?K"1� Z���aM8I8B��W��eA��`/���#+�1^ 4t5V�&��w��K�����}���|XF:A?��9���!4z��v���Θ��'
��D���. ��ND`I�zѐc�x�2�:�OWʙ�(��i�۪6�tj'���O��_E4�K#��8�,y֔��#ϐ�+0(�@0��>�����^�`?�N�"�,^N§�`C�V.7�d	����tO��投�LYfBYF�e�c!tM�ֶ��:���<�O��0H��q~��D�����j&ԧ�n��2 n�GB���k�0�S�0�S�5�m��� Ki�J�>�ʌoQ8��b����.�7�ӧ�~o��@P^��+f`�S��񹘷� :���0қ��04 t��&c��L�8Ӧj��`
���D6,c;��l��xv�������X�Ϯy�{��Z�	|s��c�c��5X��*<��a,��O>��}�i<�ؓXl�����`�Ï3��8g>f���|Λ��Zv��Kn�f��\����|�����)6O;��"̚���I05����L���&�΁���z�r�l�k	�/|�Vv�n`;�rlv�@h�<��s�fj��Zc�_~'t@?�Vܞ�z�G�н�_�}؃o1�<}��"y�ϣ<=�ϩ[��o8z±���	��n
B����D� �Ξ����5�P�TlHp��XG8$y�i~��y?��#V��3�/'��öI����H�;ր?�r �M��*�z4mi$�е����</3��ND����N�6�[����/y�K��ҥ�Oˬ��s4�.��H0�Hc��h������`V����޷3��j��5o�����Х��`�O��&��t*lX�sy��)���xc2�ݘ7*#�(�Zb�W��H6E���0�\��&�[��`oud;Lx3�6��l_<�)�@�U�B���K�Ȭ)5�^]^��gؔv�q0�A���9����`�?��`Jׂ�i�����6��-���~Z�c��x�c��4�m�1���guxS3hI�o\�,oD �g�:���mRoJM1�9� }��4��F���ɬcj�V�N`�Sx��N�FM�q���ئ(L�Mr2�R��3�P&rܴ9~S?�7��o��	<i�L���h�m`hȴ��	�ț'0^e�t��h�5�����$}������`j�,̐�f|*zܯI-l���8������Gt�u�%X�,$	��K�B�O֣ �<?��ఛ���N���4hl��Ql�$5�飩��������t�`�h�K�C8F�Đ�/�L�����r������lg$�W�ֶ$�H�g��cx�F��	$+�$���9)�,)�!��(���H��$�y|d�a���$��1JM���6��ϔ�)깦q�ۓ�`��y&j#0E}�����,͕��X��Mf��Kfj�K���sAf3;j"�I�Il/Y:��'�ŵ<�|�Si\�g��Ϝ�j�)�ŋ���o��	��,�Z�������l���e^%��Q���Pu?�HT�]�I^�#��2WYB���j@ ���ږ�J>���%�R^�'�V�S�W�Q��h�M�8B�B�h @dGi1}� c{���4�O�>N����9��q��S{�/-(tPx�>��|���风	��|�g_3��4���	��`���r>�Wg���v:j�R��v�S#��G�h-#y$,e����3R��~��z;�#�v��_�J S�2�372��!ɫ��%m�}n�!���[ܡ�L�����L5i�_�{�u/>ۉؾ����M�:@�ߢ����u{���o�F��(^/c;�`)#�G����W��X͌t�3#�k�,�%�#y�&�(��kpG��z��D�����W��ҿ~-Q�������	��b �L���W�)�]�  �%��PYJ;��C��c8�R͞
\H��dY,%�j�w��N���䓷�ʳ�ShL��ؖ�aLA ��`
�A�,c��0"��	?�{x�#��̩ �Dy�T~r����|5�:�<�	�Z{�1�u�Z��A/c`�K�2�GmĘ8'�؀�A/�w�t�Y��._�Q�Q����#dy^�V���#|A���_q�^W�X�����Tg�p��lW��t�4B��,� ��3�Ϥz�BJ��?c(�"���~n"�:�H�8�	~�� l�1^�i7���Ֆ�*ຑ�َ�r���2Vߪhx�u����nOx�"�L~4�L���E\u�	���9v�<F˧b�K3�i�|KC���r����t`�5l���x~���e���)Z��@T�tm����aAV^V�L��3��m��'|*?㝋����F�@�k�[y��K����Z~�^��
_���=�s,��PhM�Р�H�G#�4��K���a����W����Y��Jy3/�>��G�Ĝusa��?��?�˖��;+�43���$L�c]��X&l<#�ĸ�C1~�hi����q�FX��1ż%�X��,xx>�?� +V����H$���/"O��,�=��E����[o!/+�^�ϧ���G��Ï4����V�y�\��Sx���k7zzV�����6K0s�R��̔e��%�V3�F���x>l���⋎06�g?g`�t§�z+��s��뙇��a���]��-ǂ%��~��س�ի��q3���̌1|�D�4=��%|vG���[�?���0l��<3�y=�e^�a��2����*�<�	�N2*�*�Y o�u�\���% �J7���|Y�	2������x����{�����Hpww���!$F����p���}������UO&��{�����u_�]�]]]Ow��e���	D�*��F̶�ks���߁�y|~�h��u�#t��#`��G�/����jʋy�%�
���X�J��Khʆ�l����'��ՇP|rB/���V��(S *�9Z������ݮ�����F���4�B��@��RZ�Ս�N���-p4N����C#s0��q��.��^���|�������+_�����b_�ƒ���xm]���+U�G�ց���\n�f�0���l۲!!b1�h�k�A�8��`�r4S��:�xIw��K	!h�/�!��|)vsN�s��/o�ף:�zu'���`�"�&��<��i�1�P�����T��}3eb>�rٕj�'4��y�� L��ل�E+��z,�}9�^��>/T����
�U��'���R\nl+�6�}!|ޅ2����	�2o��?�p�3ϕb2�1��y�FZG�G�c%� ����6��u�3x�c�a�'��1b���mСT�u*:��'�?B}ىLK�@�O8����}z��KC����q4���e "��dt�N���F���l����Iz�#�l �ЅK�I�����d����1�Mp�Fy(!{[�9П�l������)�s��p�������Ψ�Wh�7S����5`4b�i�X��7'�iT��3%�j�M3>Ǧ4~��F[s���W���6�2#O6�F'�%�gƼ�����R�E�|��^�'`l�u�R;�8��T<�\��MY���xLL��4�d]ҵ!l,�x����=؊�����[�[y��o�kUX��1,��8���X�����hЉ��J�0��{$��c��lYG��*�&�ۀ�P�ּ�N�7;JB�;���I����x-��ݠ<�:���4Ve���vm�n�R�K���JX�
5��Ք�T�9���I<���k"�(vpm&�X�Ń)���Y���*o������ʺ��F�,���>�,�)�(�K�T��om'~sm�������f3Iy;� ¥9���	�)T�-�ؚ��XL����9�7h�>e)��SkW�a%��i�����' a�g��T	(5a��Ly=>��4c�Y��o.����q�m��Z*�VڲX�<X�g����9k.y���c+ ��S(���c%�g$�٬�"���	�@��|�����~��w�O�5�k5z'�o2��&�I �%�\F�o�v��2 p6J���L���7��ڍ�f�]�(���Y`��Y�)�|�4��)��?�l'�K�̃����"k~W�Nf���4����;�0���r0�h�)	�� x��e(�I��^	����2���#5����~���X�'��&�� !T<���d�Ӎmt�Ҽ,V�a�-E�Pt�E�� tN�À��)�B�|�`~ l�уv�5��Nl�{�CWB��^�v��/�Pᮻ�1dc�m�Ɯ��p$D�[��y�1��W�����	����CWBP7�V��	Q�����_�����/<��3�ݍ	9a�ϲ�	�`�7�j} zUb��,ݑ�e[���å*7��ʋI�xT}A� ����B�ƦK��QX��y:�}>=_��gc���G�['��5u�H:������EZC&2�e!�.�<�3�.1�1}�8����`2����ݞ�1�y8�x�̣��3
k7��>�^FP��P�@�@�Y��O�*^�C���#�f[4�n�QP���K_PO汊e]I�]�r��E���-K��2�P"�3)|���`D�����P	��@#�:���0�ǧ�E��<d+Dα"d�G��t�nOA�N	�MC,�%j��F؞h�R��B����c�`�)��d,�/��yS1s�8̝:�'���!1�_o���]�lake	+3�Z[����l,akc{{t�j������Dx;i��h���X��U~�X�n-�W���j�_�������[����^�Z���D�E`ɂ�p�1S���1r�P�.u�j���4~2��Ip��8
�4%�2� :',ĔɎ;f����+
;w�:�5%����s'N���c	�#&`�ј4i�Nu��)s���������ѳ� L�>�V��b7g�8��{���i#��G��m���J���ڵ��9��0d	�ƺ`^�b�f�DԮx�@e(Ѐ�|�w�����@�	�>[��n����@��oc�ϯGѩ��&�V��P^P/~SVf����+����ŪR?x��be�@WV�`�����#�" 	U��]��˷���Σ��fD]��[�1��8��O�s��N�J�H<�ʻICI4��O�%��1$�9���� �1܋KR�C9���B�<��;���)l��&�|q����O΢��s���"�?:��w�"����|���;��w!�Ib^��v*�>څ�'{��E��Hx�i�@��GQ��I�}x�T������>��^��'����*�:�ʯ�3�C�{uR�#뭃�|� 2�܏|����?�b��7Q��	$F�F���|܀�7����(ey�9��7 ���=�C�^��9~r��Cʓ�Hz����<O�/��c�����Ox���#�1���!�wU�_Ćo���+(���v���G�s"_�}��^����C,˔�|�?8��'�tw_ކ���#���ن8�������"^�o����Xq��dǓyp�T�5XA q'x�Vr��z�ڷ�|��R���	�	�K	F	Is��/�q�HC{!�4��f�-TӹL#@ʔ.S�����2��D�s�q�`�>�c	�Sȓ���\��/c�1���t6�Se$��eM8Fp�{(�`��nlP��3`א�.��v=R�����w�M��l�ڎ����Q���64�e~���~dP
	�5�%��xF���%}�dt��V3�ρ��{���o1��\~4��nY�=���f�;��τ���.e.�:���uܤ
v\vb�[�����c���-d�_{3)� (��&b�1O{�JH��i)z�ݗ)�e��n��>��{�w�E��~� ]	�i�)�Õ�iJ�4�L� j�2j<ZK���4��T��oQ'�j�4m��-g�V��-�8s�u��5��^|���XJ�����h<��B�x�.�i�Xe[y�x=9O�m�*�j���=����%�T@���A��)��}�o%��ͱ�&�j����*�,U�-����D���.y?ͥ ��ī� ��i& J�^%�p)iψ�)�Ѧ����&͂(����OM8?�E5��m��ψ<�����2�l&c^�H=�j۔�5?���y���cc�����w�ǚ�QK@����������3�����l6/�|����R�d��r�e�cd��7�WD�v���l.C¢,��粡6zg2�tO�2Ժ��	���jQ*��`������/]��D&�	�&���JF��V�N�l.��SSB�l�oI£�3O�I��hP�����+%_=D�oc��rXׄ��h���+�N���TX�K���dXd��&��p3vO.��*�C}1f�/A�-�Ý	*,�N�Na׭6��>{)�/�#��D_;���'�q�$��D܉lz�j?yo܁��jB��*���$t=,������|86�Rѝm�A�4u�N��|�������~�W~�W������&P�E���q =R�a�΄�.�΄A�ĕ�U�ӟ�����P��2�����`�)
�}�: &U�`F#�[�:LX���ȹ*�����a�y@���@A��x6h�v�Ϳ&�"�<���OH��4�	y��&�8e:�³ l�$��G�jT\ڀx�k`i \�1�s2���q��j }¦��hg�t:�������0�m<���#�x)�|}xj�[B�j��*�E��7��+	���U���
�m���,� �Qt�. �g*�X4��L�MW}@e�O	��GxC�#�o� P�!�t2��!ao:R�e"�Hr!eo6�����!�.���$��S�3h7� �Q��"aƚ���2��O%�����C0s��O�fN#Ѝŀ�}ѳG7�w�E�n]ѭkt�����ll�ѹ�=��:H�a�e�^=0`� ?é	�'�a�9-���/Y�c���P��[`��X��{�s�6,wv�gaִ�<~F�ŎX�
�'N���s0k�"L�>3f,P#��趓&�羅�Ř5�I<4o�;""2�|��]���]1w�3���)S�2m>��[�Q�&�r�����i�;F���^}�7!x�ԩprw�J���s�c��t�}3St��E���T�K��M����c��",O���G,Iv�;��=	������ ��� �P�-��� ����u��<�'�UP���]W����g��-�˳��Q�%밲�+	�++���ʛ ��"��R2Qti0RK�p���p�&��D".o�2�Sǐ�S���HB�pjӆ��B�.E�wZ��T?A}i���%�L���SLq1�L!��ߤ{ujN��O��8����wP���|cv�v�s۹��q6<ڍJ�a僝�zX�
�g��Q���Β�Q"ˇ�܎�G;��j�����b�{���T��뙗lo~�nBh�+�w�+[Ptg*���f^w+t#AwS���L;�=��m|}�f��,�����w�Y���ZB�f� �<浨��<v3�o����&0ּ�r�݅*�x5Ar�]�����Z�x'����__š�/����������܅һ;Q|��\ޫE1A��`\��~l%����6}|�,o(#�=أTC����y�����p������aˇ'���\AX���)l��Z�||??��_�Ŧ�Ϡ�X��I�_�+	������G��ro�Y���WY�zm72�Q��|���"�a�_�CA:�F�ܟ��$<�G��;|c3Bnn!d��w#���z��G���L�<omê�[���V8�ۀE�7`�j��]��30dsF��T��!;�0t[*�nN�ЍI�_�^�ca�ϒy[6�]O�ץR���|:��S�+Y�1��fF��b��˘�FhH���t��Ӆl�-F��S!ƞ~�}Q�ɗƠ�b�)c�Ѱ�sĀ�&�H�9������I�)�ς�5�T��}��&a�,�xleiL���,	��<�V��W��]�
�8���|���`�`��n�}�@�EW�q'b�� jI)m�g���}F�^����7�9��\WxM	�G���d;�������`�=W���F���R�ym��\E("�W��d#^;��	�q] LR��c��<%^O�n��	�6��?ds)���9M�e���A��lڷR�ձ��6MyVZ)U�T�Rf˫)�ƫ�0+�$맩��ZP-�>#	���0k��B�,���}�j�G�=�,��b�:5gyd�x-�='����9F,�1�"2��Ӓ�8o@ �绪�gK�h32݀2`1M�K�5����ϋ���B�T�xK��oj)��3�wD@O�'
B%]�嵛K��@�o�7�-���*�X
T6�����G�0u	���������T�Z�4�_���'X6W��i�x"M��J4���xF��1M ��)��t��2& 6� ��qxӠ7:��#ԁd��0��M�뙭�z���7\��X��]��ՠ?r��59�
+��%!T�r����@4�x��)���=n�G�}���oc<�5d���<tݑ�t/�A������x�k��?��S��?~�����	�S��w�}rK6�w�?������$t?�۽)�"�d�EЭ���̯�@�+��	�d���������y}�m��)�
}̴󟼍���_I��\�n5�)�	�b��o�A��'�|��û1*�ݳ}`W�*�@5)�D�boL���ӎ45ѲJ�P��E3Q!"dd[��[b4!�� ����d���!����d=�  �Jٛ�ߐ��S%(<]��}Y�c���X�,�Y�����wNo�O��A����/2�e�^2'xZ��vma�C�}Ma��f}L0�u22v�!�p)|	�>�ch��c��(��s��e ����R+X>��
�4e���=��|��4(��[v'���	G��$};	�	|~%W��j���@����YO(8˺=Y����H�KE���(GΡ"��� �.�`.��d��MF���Ep���U��-�޳0�y
�,��)S�b�a�>v&���ԔIh�0�7~��}��G�^������%��l`cekk�X��κ�������vB��]0t�`5=˼��`&M�cL�8ә��0��<�9pY��%�X�ꂅ��a��b̝3��9��y.XW,uZ�Y�`��
8�uĈ��0~���D ] �t��Yj�iS	����X�lV�X��u��L����RT`�ȉ<h�_��K\1t�t���ǌ��ŋ���P��6y*����������o�v^B��Bk��nx'��t�{�J̋Z���K�]�8�����3�)��<�{ �6��YR}@%W T���iX��f �<
k�^y�O�5�nY ]Y����(#|VxýR��z�c� h\E8���q���x���(8��W7b	̩̱���Q\��Y���V�q��;���ɾfFcX4��ǃi\�a<�b����;�(�ץ��}t�>��-��۵��#���W6���/�V�ҫ�(�\�<�yl<s�X���2�K!a7�V6����l6ZeҐɤ�����yn�ʻ�chtg��C.�+%(�u
XFY/�1��΢a�K#;�J)�/!��z�����E��"�3��zJnV!�|>��B�E4�sy|��BҐ/�V��g��G��<�Ө�:_���5Y���ը���kx��(��m��\	�.Wb�-�J ���Vu\ٍ�RW*�s�y3�����b���j��77���F��Y�V�E���J��*��J������p�>!���w�w�)���ۊ2£�}���T�j�f%U�p'��P*{u;�_ތ|�5�j%�y�"����f�o�n0��;QE�^�j=A|6?����a׻'p�+8��˨��<�d��P��al��v1m�簃��>��'�P��Q�b3��B�k�Q����yU��@�;����
r�]B��x�j޽��，���w^��7o��X}d#��l��s�`_�·�Ї�i_��]��>���Ԗ��1���jIY\ʅ�ŜeF�49�I#)��Ps�1�+C[�4e^&4M�ї��VB-P�n��XY� K�*^@��;*#[�$lJ����O"tj�4:Yn>�f\7罘�~��L��^v��ښ�h�gY�����P_k���k	u��!�*�vH�H;�W�	��wJ9�A����I3I8�������ߴ�0�X�r���
%��(�<n�0���ƵVO�jܧBH�=V Z�/�mR	I��c�9R���4Ws��_�c[�XLY�~-|�WW��5�_A�xN�K��Ae�i��*�X)�B�ấ>��y/M��hK2�%������&��<�O M�.O����)�a��iT��M����_��o&�����d��*Rp�\���8�N=���|OE�rn3�s����}�uV���D�xʚF<h%�����-OnӴ�M�=�Z�t���S@�K�gmzK�&�$�&���OJ�O�=����k�\z�^ͦ�Hu8C�<���Ω4�;���L���[�i�s���'[� �H����xA���*	�jA��D�;jx$�9	8
�
x���ԡ��t6�H�ޮޕ�C�Z_Q����;+0~C
���)ϧ�kLഢ�(ɔ-��q0)@Е}x��}��o
_��{�،Q�	R����	�p�g�}��~�	��^O��SMs��ݟ*ؓ����~�)n~�>�|�.r.���8��D	�CN�W}:�K��3}�n��=�����k�����_��#���gn�N�ƽ��+I��G����G�y�I�a0�r�]�7l�ܱ�*7��H�����_ �`-��{�.u5l��`^�#�F�kХ��GÙu�dc�S �A�d�Խy����j\�,|:ŋ�m�MO��`�)�wU����O�/���֕��d��x�%�a��Z�V��Ю�Kx���@����ſ�ֺ5��:<;��Nf]�a��v��a�����c��YH�I�n	�@H$�
@J�����J�m�B�)L#P�ԭ�p�
W�_I�rW�\�M�P�~��ޭ�ӵH?�m���x�f2�g"�H&⎤#�ϬH�b	�'��	S �?�u?Bh��,���w�6�R���D����@ƾ|$��D�LA�#��I�ޗD���h�[V��o��lLw��is&) �  :n4!tF�>�z�߀�=v4�O��q&&G�����ҵll�����]`k�	����]�Ӿ�u�##=XY��[7{�cƎ 4N'0���y�1����k�V����f�PZ�hV�tGLL��2W�_�d1�������.��X��n��g����cX�6��9�����ф�iK�T,����	����� Dr܌������5�0�@ڧ�`�����w ���}����5�0���վ����%N�3|�:w�����ڡ��齠��1�}*��ݱ �K���SF�ݓ���D�@` ��� �>[DA*we�Z�����H����>��A����"�.jеX��׽��K�r��++<[��|�@%�`��/ㅳ2
������w�c��*��F* �nTa%^�A��1�N�%r����Fe�alTG���9=GGР�I�G��q:#�b�,<^��+�(zx�?��K_���W��7��B6�Ji@�P�4�
4�`f��f��F4��b�-�4z�h�f��U"hJZ6��,�+i4����yȢq�y64�E�gsTZ��d_��,���PJe��v&�����iܗ��6S��k�5yN&�,��4�5y�(�5�N�\*� ��cDi<&M�)��\�S����<�����gy�g���\�gb���Z\f2e�P+��D	��<q.��|ә�.e���Je3M$�,k��_"��H���~ϗ��^XO��,�S:�%]�d_�T֥�W�"��d����ԉԍ�/yg��xO�,s��8˛+`�gP�|���zl��;^�C�ۇq�ӳ8��x��>��I���.�x����_F������B��n-��~'�����-�ߔ�g�*�)~�c��_�!��}��w���{ "@ݿ���7���;X}l3��NE����{���z�a��Ȼ�y��]�+j�{��saJ02���*�iACX�fL��4+�үЊ�i��˜ϕ1)3.5a���ZA�y>�"3��9���-��h�x��h��@�vJ�x$� ��,�K���	������4�SIk�gC���H�c��t��d)�ϵd�6|�_����G�!�vb���AHCN��$�͘ƛ�%�9��b�2/e���5�	�j����:3#蘰>	�Ƭc��r�Lct,	>V�.Y��[*^KY�9�
��4�TIS^W�kʼe��"���Z�Bym����l���:�����ƛ�C~e_s����cD��-��I�uB��mͥ��_�rډ��ψ�6��*��_-W�[�>����*HmPy&dDc�x�u�!�M����z&��f��7Sޣ	�d�z���ߓ�et9� �g�i��$]�D�\7`�!�Ԉ�n����"#^א�p�@��E�O3�3^��wpl.I��+�s�ѳ�%R )��y�|?��$>��\v�q"Y��x�C	 6^O�j�1�����P$ס�Xf	qV�sY~|�:����L��2Mō�k&���:P�I��j�����W��M���xJ��	�"�WBm,�<u��N�(��z�iӕ������0��	���q�Q֏$���$t8��c<�x*�y]��Zq�EH�?��T�2��V�0:����9�Ij ���q����	ی���|�)|k+0�0]h�[Z��$��$��|K¬�xV���"�>G7�	�_������G?|������U1��19����!�c��|�������o>��?~������	�~��|��|�6۴����޷_ �~�憣s~ �lK�}Y�ɴ
[
�������6����������[8��=���5}�6�vg^�����OYF6���׿��W_��h�*20 �6ދ�RI�� ^������	��m��(ئ��U�/��}�OcU�p%��`�H8צ���e� =Z�\Qb]B$��p�]�oD#	�2��H��2L�tS4�c��/'���B��G`E�J8�s����y�l�[¨�.ZY�������he��c���μښ�E;�6�5o���5Ձ��.L;����	�Y������3I�3�\���1�aW&e�!�� ���v���F�P��f��K�S9F��
@U?�H���h�-!��\�#�{�w0���R�t,����	j����D���G�&�� �.�vj.mF����8����fl��%�*�q�п#a;���}������J�'ܲW�-��|�b��L�4��Ř��0Q q�$L$����]�uE'{{t��#G����S	f�	��ѫ� �&���1�{BW{o�}zF�^�`'}Gm�akmk��-���cG$a��ep�X������·ӊeX�Z��DPd0�����GWG��^�Ů�p]�
#ƍ��ISp��]���~BZ*9e�̘2����q��w��)s1j�T6�P=� =	��������X@̓�RW���{]0���FNĀ�cХg?t'���<k֭C|FW�ŀ��`գ+:�@��C�}k�m�"^l�?�龜QF�1̉��e�nXS��]	�$��F!����J��?��a�+
��/����T��5K�-���F�˹�6��l5�U"zK*B�b�wǯ$k�ᚾN�p�\���(�%�6z@@	�
@��	���XK����p5�J�!Q�M���g�wϢ��6���³Ř~�c�Tc5��1�fF__�ת1�0:�J��S����0�rF\�$`f`�Te0���8�N�`�<L��vNb�,:\��G�q��O.&�
u���h��G�Ps�U�r��@g�L6��lS�p��!K>��d6<)l�Rh�6�;�H��s)J<Η�@�	�d[{����Yj_��S"�$^O�T]_];��Ee�.�$�u��Fx4?��ӑp*�"6h�ܟN���B� ����q���8ֱl�� h�T�����0�$^C�H!��e�)B5�%��W
�d6�Z�0M��Ө�N�}��~������N�a,qG{$Qՙ�W2�P�.���-���~�-��1�4�h�D�H�C�M�ke�����F\��^��.}}�^ހ��*P{+^߅=w`ǽM� ���La{d��h�)駊P~y��y�~|���wlp��ȿ��·���������_L��WY����c.��%R��Ɛ�$t;��F>�U�s%�v��N���|��7���E�#cޣ	�O�łF����F�l[�X����-�D8Gԙ�gM��"�	Tt"\X�\>	���!e�H��2��v)�Q#e���RH(�&����:��8�L�kL���U1R_3^[B!����ƀ �6S�i��Ĉ��ɉt���m��w0���|{=dTdK�c�P/���ԅ �����4P�g�Ld����NX�bT���4�sΦ+ɺȘy�^�5�	OV�(	��pP	5�k0OI3'�hCF5!�b�f/�����	U�"�W��e`��}lĠ׷��Z.��u� ������ *@�I@���,� ��5��W�~2�p>��K���l�/����#���_!t^�h�T��k/�O��<�M$5���6��z�18�d=	0�3�_�H���uO�G�H�-��k)�5�q_s��7����M$̎|Ve)��Ji��R�)Ϙ��]�mY�ȼ�K��l�ť@��'ϩ�5��9V���k�:)/sKR�v�
��p[��"ޓ�ªP\��ᣀ�Yi�s�ג���ܣ��kPY��)p�LڐZ��(��&�I��;�s<�Jj����%�u8IhU�'��1�ڲ=�p�=Ձ�AGV.u	��Vu8���+�J��e���o	|"PK�١DX7$��2�*cq��7�)���+_��=蛳=h�w�&,��8K�9�`}4V��`��+v��߿Ə���7������^��%���ۍ[�|D��_��z�p��%�q�o���G���Cι��>�u�_�k�}�/�3>��|���x��Whx�>�D�K�7���A��wq�����O��	_��>��y�b�Wb��t,"�.ƌ48��/�#ز�����o�����~���~��d�-��y�8��{��f�7>�y�v`D4y9L�=ѱj:V��n���Vb��8mO"|E��p�%�GJ�G�8�>!���͡�L𤱽1a�c�;	�R��7��s	R�X�G"� �.�����;�������^��C�w��k�:f/��E+�Y�@�H�F)�7lC���A�X�u`�����a=�����8�I��@R}6���^≕���D��p���R�k���R� T�qUX�� *Ǌ���*��ՍϧxV5i�H��WS����Uh�NC��D�C��Î`.ÑF�3�0�n} �@�Ԡ��T�ި���.�ީC���9V��~F�CԞ8D��v��EPY^�Ar�K�<f`��A1�7&����c옡�3g:&M�aÇ�7��O��;`0z�����b�)3fF�����8@�sǣW�Q�ҙ�u���F�k��066���;������076F׮�5~0�̭����f:9`��9��S��8�I3k<FN��SGaӖy�c��,w��%�4z9",��� ��e���J�r]_�dHh4\��V�
��2����c�p��%`�"7L�1���5~�pX�A#&�g�Q>vFM�E����3���!�p
����`?��lM�c@ m�۶A�v��k��¢���[��XY���q�oHU�4�����%tr=pg$Bw� �!A��H��' ���t<��`M����.Gޱr�nMCp�
�_�Յ~X��%)�p�^��E�X%����^�����oO��Y��POB�o��J�^���1ȮN��kG�����Pvv+��U��bf�h'�� t��
�Z��J�^��4 ����xe�l�7!���&���A�v"��.�>ڏ�wO!�s�{��^9���QK�<�͛���Gx������}�^���(?U�R��`�<OѸΠ1�v6��C(<��861lD�������$^�R���M��Yʾ$B�6\A���w���kű��c�4)C��SI4�SX.-�6��lK�<������p��,�f�L�#��D�qB��2�0�g�t%^��E�_/���>Q<̘#)�^���Ȳ'��/��dWYj'��4Y*�d�s8AAf<! ��u��m�߿	U_�k�*��4��X��9`�h�0�h1�yͽ1( ��?م#��ǵ�e]&6�"�>quш��VɏmȮ`�����@�h���G�e��F�@)��Ǎwn��?��?~B}�~��~���^F��Y�}C}@P}_!��3U��އS5�����L>��.@ϳ����a���W&4�Li�YР�$tYиӮKI�o��r옗�����0�P��f�>%�R�V
����3�!)S���n4��@�d*�/s�u�Y� T O�΀�����a�*[�4��2P@YF1BŨ� �
.e[��IX�>��c~z��Ӏ�lDY��Ӄ�n��7�0��Cv��
�;%S����>�����EB����m)�W}deI�5a��x�%�7=�WS�d6Υ��@�s��O�5�$L�1�4�5�p5בm�(�>�)��ڋ�6%��u��jw�Ty8m	L=�V����>	YvK{Bc��%��o�=e�L��׋���������)�U��"��tK���\2�;NJ�(�4!�J2�TA��霪O�� �����\j�¦@U_eޯ	˨�O-T�9�G��ϊ�)b��7P�@ᆿ�Bl
ĩt^[yI��!S�g�%��K��sK *��\O����T�C9��l.�h�@�*7���<��$��c��5/�x>[P�zs�{������G�Z*`l�-I��<G�O����K��PQr<�@ū�\�җS�B��g{���;�Rj]�S��6G���H�	�R
B������#ۓTG-����J�Q�l�(C��"#ʘm��xS�q�P�Ą�x��u|���ɟ���������2}�{���)�kp4F,�)�o) �;�ri�՗��_�K�맿��7~d;s`'F�����D���!��Ox���k?}�����{%�vbEY�bz��d����UE����_�a��=>��{����.֫�6~�1�,�zC���e��O���Ǹ��C�ۃ�9���v��+i9z�8�w�b�T<6�;�[o?��_~��%W}7���9���S<R�D_��+���s�u{16���n0)Y݊��X��<Wt-X��#�-n5�p)���D$.A��*��ޙ?B[��D�C\}rN��T)R	��>�o8�9c��l�[4Vc���G�l_Ŀ_��/��F���m�^BG���`�:&/������%虶C��hO	�v���z�:�3 |�E{c���}�`7���a��h���E�dxV�bu5�!\��
X��i`S����QMW�6�]�)��`D-��zn�P$�Pٿ�y���	�)G��x�v�>�j|>#�RJ{(q�=L��:��MW�a���(?QC�G���(<V������Z�6���� 	����E�����Q�0�u�M���cЀ:�/ƌ��ӧbذa2t(������1�4Ga�C0A �QeG��J �y9��>��J�N̞���ݠ�kks;�X�܈21���!L,еo'�0S�O�T����yS1u��"��Z�I�*0u]�k��a��+�t�r_o,Z�)s��U�Ќ�\�G�(�\������k1m�|�;}h	��Y~pt����x)\Wy�}�?F�����apt��"B�%nX���T���c���=��m�cH �!���s��m۠׸>X�Uy�pNw�
�h$���y�m��'��A;7�vnA4Q�ģ���`�_+��05�
ť�Cr}7�~��� 4`S0r����ĝY���e��-	�� tM�Zʋ���rox�y!��Q�!
@3+�����G���9_�˕�yg�@GS#o��#/U`��r��^��4~y�ߣZ�|z����m�^��//b������m�}q�\��w�a�[g���)4�}'>��k��=��}���4���_>ı[{Q�/���6��p�l��&��D1/8Ql8�ī�t�nIQx�3r""�%(E��?�NYj�K^Ij_SI��*�/�j%�"�B^�@l3	X&
7��o�3��a��U	����t ��N9���O��l�8��e�4]�h%p��/����(�
Q�x��c�nK߀�}q����e��_x}4���:�:���hDpu ��Z?��C̯N#��H��D7��:�ԩ�lA
8�3��F�H�:�x�+vo4_�4d�H������,_t�sw�e8_�`��Ě-����²��������#�9e��%9y8��4~-!H���w~��)�=����\~���F��j������F�z�(�A�z:�Ne��+�lN%��X<�h����3,�L�i#"ĩ�D��$%�&eP��ҷ�F%��ݮ���
��7��LvNRM�4c~�P���<�y��*2��A�d4Q�GdL�S�Tţ�OCP<��4�%�Ԕ���T�S�'P1B���=�A)�{Fh��>u	���=��ј@O�.3=�3�yԓ]�p;z��CAh)��"}F%L��p�:֔�%�V^�F��K��H���z�R��j����~��W�h�5	�"=���,O�uC��i̋�W���S ]��ȗsD��&'���J�^S�͂�Y��N<׎�g�|�X��W
	�E�|�y�LxU���Mƫ!P+;�`gh��|.����=U�Z+�!��!"@	�Z ����TH-�>EZOgSiAT�� �������I��p# )�������0(�ƺ���СQrm��{�WTA�U�ׂt���=/��j�O��RP�**���)xj�)�FO��Q��f�fK �ұO��\���@����H*� �?�l7�� I	|J=PO��M�����5^K$`�\��)b���a����+�j���I�kC�>�� ��!P�m�ۓ����o�H`T��������}�ʀv�!�J3�a�6���b���x���1����o��y��U� [�f��1�h�2��l�l]
i��-ŭ_?W�����wx�×�?���ݱ�8	�~ք�J��ß�����¾�."`w�dya@���F��5�I#�G��/D��J��8�7~���/5�@r���	p�̌ �|��~��?�ş?���K��Y�Ņ�㋡��D��5
�	?�
|�)vl��#bO�|��*�t]y�o�!]�gcR���uW�$�������P}f?�Ʈ�M�3�J=aXN-^�W�,Z�難��m�[U�+�	L�:E�<S�����!���@ɹ2��C<4R�)������?l�Z�m϶x�k+���_���i��e�ښ�Q�h��t�:hg��Z��~+�p���5:��t�����L�`h�u=��nkt�oM m� �j�-�L��s�a���X���[㱶2��52�J��M~��2���۲�M�5�h��	m@W	�J:ӔG����p�M8�����%i�E ��3)6ܞBhף�F�E>�}���z�V��x@+N�GFC.B7F!��
`�A["���%�D6�cݖ`x�2r�by�k�L[0S��Ÿ�#0f�p�5�@9����mX���`Ĩ�4x,�O�M@�̩9��6z�,̜�77?L�����ǜ9.8z�<b��ѣ� X�u��a'X�u&�ڨ�,�	��������&��4���4{��F�-�������g�򃛨ؽK�<�x�;�,sĈI1q�,x�b�ƭHK�A���v��Zxx��i��V�y�&M[���&�ߐ	4j����qS�c�>�3`����0m!�Sf:c�lg�=u�#Vz :%��)��G��oW�wD��|6u����%�a7�3C��<�Cy@W� �.�g��{Җ'`J�7��sk ��P���H?�9�>��#	���m�7AU��	�[�TBp}k��u��Ф���� ZN UKBh��L@�/"+��\��$\�u/�~�4����?U�e�r�nU�A�@GP�n�Ǩ�L�V�I7����xk?r??���a����������!�z�8��9�]��`���}�����q���q瓇x����ڧ��D�����m�����I��t�):zB<g�A#�R⹌���� R`I���CK�������7�|I'����������Qm��h�C��OJ��ȋ'	���J�=�!@� �mTܾD$�KB�~���0*׌n�(�EI�y���ͯ	H��5���:
�B�"Y����#8�Ux}����=Q��h��R�C�0�KZ�/� *@J�e���R��*��7��p�7����,O�vI�QQ2���P6|����#���khm�E#��E���_0�'s"�����J,�����
�4��%�[��=�/s"�N�aϭ�8��>�N�}'_;�/���'�����p۟�y'21�t:z�ICO}]hxu!w�aՉi�'�`q<�*�+dE@�~�2b����"!��$���r�>W���R	�\(D�K�.�O�Bs����M�Gi��,�2�Ȋ��BE�.ǘ	����B��;J�Y�QJ����(��wM�T;_��P�l�a�{�m�bFyT�F� ��g��L�t��5$��x�m���
�{^/W:蕍�V&�۠�T���|v-YW�̻�$?	Y�>�2hN߇[Ԁ:��XƋ��aǔ�Q����Z��4���2��e�xF	�<K���*�'��c*�)���OCJ�y�riʥ"e�s�	Kք%�?4�u֧@���=�ѮQ�ޅpו���JA�=��7��Z)�ez�����r�(� ���j��v��μfW�� K ��>��Þ�����/so��ɜ�j��FYRπw����5�a>+�?5����YD�S#���z>���)�lE h{>w:��vg2���L��VI��=�3��k.B�sb~-��^s	x��y(I_\���Zp�P\�Y;bkS��{�����c�|@e[қK�*��T�[�)��� �
�m&�Nx�4��O� �ߠ*�����,�I<�ھ�Rm��+�jBn�^Ͽ��ա8���p�����=��l�t�� �F�?U�F��(}�i"ʐ2�%�)�}�8h�?z�����7���#�c1�$=w�8B�)�'�i�2��)�6��фF_,�]�K߼�<���3��
N�cb��N���{�ܧ��۟��J��wM*f��aXy �nCw�����ѓ�_�]��U�~I���
{?��'�����>}�����;x	f��a���?>��_���c�05jǭ��� ���[Ca�1]7�����A۠Y���;Gp���Q��-�]l���0tZ5S�|p�;������_�ɏ�`��Ø��a�*��U�/X�,�+�Ƭ-1X�).ap.	V �wv
NW!yo"��&!�U�cn�|��ٝa0L���/vz�:���{��[�}W�ضA+��C�|�ۣ�It4툎\v0jO��!��@ϰ�F:�5h� ��ް1W��@	��5� ���.�1�7���>�=s-�w��gCVׄ* �t!`�4��	�u�P �W����COG�m@8�6���e-ω�OD��B��A��4�v&%6�r"@w<���uK�'�>Uy;%��h%���'�u���MVa��;i�G4m��}ɴT���J?x��cI�R��;�&Ĥ�c�0gfL�N ��#Fb�Б�8y&,v�|��I�1`�8%�M�� �����d4}�����1v�\�3��MD�	�k1m�#���k,Ĩ�3ѯ�ht��C����ֶ���ٚ�;�gb��p[�%�K0�y>�/��y�!89E[*����k���K׬�1Ky�r�����u~X��^��5k�����,��Y�1u�"�`����T�aS�w�d�����1v2�a�|�pX�	S�0d�F�_��#f��Љ�p�
DpR*��xb��	���&�7�G�����Vz/�����·g�/�e+Y���1H�-�'N��I�!PҮ�A��q$�d����*�g[(!5^�Ky6.����_��
O5@U�	��q�3��G��!�k+E^j "Oʧܛyx!��)5�
@��8A }�4�U( ]z�B�@�XB���5.zs=�>�_)Ǆ�UX�`��;���Ρ�ͽ��v�˛�h��77c㝝��J�����''qὋ���<��>�|��	�����7���'����(9��\�\6�Y�F�U����'4᫲-�M-<
T�����ds Ղi�/� e�ږ}Z�@5���ʫH)�c�,e[�}Ծ�M�s���ɹ~+��@01l�B��OB�&��&l6U$��`N����r�HY�$���q��06����J�� T�8��˿FI?J�p���G����yi��o��zm�[h~3���\!�7H R��u�L�c=D�,�A�dz<�-�/[�Bi]4���c�k��y�,�X�Rw̫X��ի��f�6x�m�Vl�%���w_­��F�� �|9�qg��Bݕ-�vy��ۉ��������c��$t=�.4��iL��p��aey*V'�aMc��D�3a}��t&v�K��J��z�@"�v���y��/���y��i]� }�kx��<׆�%X�7T&P�I��(��S&Y7�~�d]��	������D�|dP�@����_i�����21����qP=��.@�K���T��J��@�@ÿA��	�KQƤxY%o=	���gF�F��y�6�i[և�ۄ7�0���zg�O��6�"�F�ZF4re��֫�\�Ш4 ��_��|�e �R���L
ڝJRi�Yn���x5Ϧ��7��4 ʲJ���v:�Ӏi�]U��)�jAY5�B	��D��z�,&�O�q�5�z� }/`��"�\��1�;[�Y�n.|PǇ�1�存}c=��(��[�~�
S�Tc�*�S����W��O�k	zȻ(��d$^�BX� p����\Pפ/,���% �T�a��xyX	��l��lY��SsO��R�M N �-��O�7�{��/�\�ו>�ͯ#�<�3��$�Y�#�*�{V�F��o*�ڐ���S#�	!ϭ�[Fn����g5)OS	X>�M���T�0�Qy)��H�� K��{�z,�J�m$É�E5ߞ�����Ф7���~���Ԓ4Y���j�S�n����`�Z
��U�~����v
B45 ��P�R�#��Rz�E��)�+�[����8�����(������m�L(�B��	��iB�4dY��E`c�Զ>�J	!{�p�wT(�Lu���Pp� �'��!->y?��>��[�z��؁���!�"a�+f�a�8E(�6ac0ӑ��'u%��!��v�;T�]���1��05�[^>��yU	�����Pvn/�%�`D�l:6���ngl6�fC �f[���Ű�rD�w�" $x``�J�{���,?y�6s���7|��w��r��`� ��n0�[	�7�e�b tΖXh����0����D䞮A��
էӏ@�0f���&xi@+�����2���uо�K��с҅qOC�u���K�h�miЫ>vT{����^{�^K��%xvd�A��muu�F��tl�6�_R!���m�k��i���n�2�;���A�#���1{��+m��
���:��H`T��si��PϝqX�#��F)/��Z�"��\��T�ʥ�0�7I�z�u��G3h�j"����j�8�}$}@öG"vW"r<��Y������ڟ��C��<��T*a?�t_���3kk��]߲ L[;�}��g�^��ٳgO8�F��(s0t�X�7���Ŕ�dN�6k	fP�\0z�,�=#G�a�x���3]��B��a�i0:w���r�,��tN���'�ζ��abd�.��1z� �5Ə����X��0¤��;b��)2iFL��\_��˼W`�*�z��T(�#��z��z��}��Z?�8��&4�ǰ�a�m l:�À����S1z�;��9�.��H��ՑX�w.��`��E
B'�p�ܥ+����@��7=��y[Y�@�c;��m��
�݌0m�L�������|"�m	����_m�v��v��L��}��	�A�Vyo���^ܨ��(.��N{nX�Bp=�}���~�RM�9���+��K �R�yU�|�%s�B5}@��!V�ˇ��y�܈ ^��b9�ݨ�d�8�稗7`̃m��S_߃��6c��RL�R��v"�]��b7JnC�[Qyj^َw�c��=8��0N�y
?��[��"x�ã��������w������/2��/nA���	sY4�e@�G�S T Oۇ�)$
�*HzVM�Rg������>��6��I(Ԇ�j�h.��8�b|3IZ�x%�G$�.��N,�y�S����kV���:���GTRQ�'B��RO��'!r~4��������aT�%��`\��a3iT��gl%n7W0�K�<���M��n.�Km���"��o$���J�&�Z��X����ERf)�����f��7@�Wcv�f:cf�f��¡��+W��f�6�����X�q�nX���AH�1�>��-+��jֿ�	UOv#��V,9��ф��G�`{,�%+�8�΂�n	O>��g�Й�j{*��,X��`������r����j�Hz]*A�3y��{D�
@	�jt]ʊ�)�)�����"����Pۉ`cC����m	:���U�I�R���#2��9ASֵ^EI��te4\M5�����~d�\P��@�T?��~��8R�%VB_	��K�Е4�2��xBU2%�ٲ������d&<ލ�lư�7a�/���t3��d:������Ret��;�	����gJ���-`�G�O��9���B��J6�/�����}"#'i2�V��5��oN�ߒ�aMHؓ��ַJ��E��]��;���]����<��]�!�K0����+�s�K	�����A|���˻�{��׷�������on�/�4���}c/\�n��k՘~�S/�1?B��J�E�j���F�n�	���WY�+Rn�����P[M_O5O+�I��$P�4�V����z5��Bv�.����j��
,
x6�x6�K�S<�Mա1o�s�^���gJ=s<�� ��J�eZ �~�υ��f�T�& �s�tx����U���6��T>��>棼�r})�M<~�2E��l.�n����R�vYʶ�uy�S�����ז�1Y*�޿\��u5�	��栨�V���.�-�{�y��R� �\/)P�Մ�M�x3���Xu�H S���B�Z��l.M� �Z��v[.uţ=P�AI`4Z#B���H�����o�DGB]�}Q��� R�!J�j\ꋱeQ8��;�Z ���q����o���@t#��)�/=�a��	��1��	�\O,ݞ����_��K�ʾ��(�p��|1+%���_��_��3}�1�N6`z^����X,��a$��A貃�)�*�`��˴e��\�^%^�M����Ѝ�Uc|���_a��㘙���~�I�1����z�A������6�`K�ո�mb�c�:�-G�Bo�.��M�#�fycߛ��?��~�۟~�w.br��.F�_t-��n�"�%;aLU0��N����XQ�奡�۔����� $���F�x�´�i�z$�����6��l��0��~0�g�ކD=�Z([�]Ǘ��JQ��Q�;t@�}{����ڡ]��hݾZ�:��Z) ��x@��"Զ�yOt���u�=5�y$�	�I�U�ګ6G��V�;,��W}=%�V�p]����S�|j�� �x;��� �ʚ���+��@�_��*�vXr/U �|1m�������&Qk!����;%�6T�/g����s[P}z
�)Oh��j���Dɹ*�*C����F\C�P���(���<�t�~f��ckkk�m�u�`׹+��sDP�7*	��-C�>#��D��$Dy�bҴE=�c'�ǘ�s	��1x�倁C�#0$q�e<gz����[GB ��g�c��?�c��1�n�c����C���&L��f��})�=�aɊ��6:&8L�X���0
\�i�+\�V�;�^!�X����X�U�>X�gg��0��CמCЩK�0�=��瀱4j:S��!"6~������������\��{v��LU���=����(L^� }'��u��0�2�s��c����ho��&a-�ӫ�^e���EFؗ�����Tv����$���99#�>��w�	��+#�j��j�_Q�m!���8
�:��>����NT"rS2J#��(��AX��|I��P�ܵXA �(�@ ]]A6WQ���C�B�]H�d���gV$�����WQzv+�.n��+U�q��h���Xh�{m&���h(����%Mxɭ��~kJ�B5����(��E�k���64<<���]��On�Χ�q��;x��]<��.�w߽�G���_���к�[��+	���Q@C[��L=%^P~|��`A| K�M�`W���F@'�NZ����ʦ�Z��n�-I�}N�k�u5i�n"؄C��gS%6����|������	d��SyO���B$#���*�KPz�%44�e
�3�=��|.մ,\�:���#He}��^��ٽ	��Ɇ/��@�x9�Ra����Q���\����E+d�rl�[ ��<�P�{�����g$�O�m�ό���\����1�p��@h(����c�Wn
���U���i�N��G�SN�^��0ꆹ��1��	.U�X�q<6{�c�/<w����Y��3�s�y���x�
.��1��ٻ>�	��}�X�N�h���s
%�Tds*VR��۟�Gw�h�;5�p;��%x����F��sdJ��S��V,�5!SBmM	r�\Zq[�p5᷹*�֜�gF𓁏d $�&���O�HF��~I12�$p�-�$$6K-�h@�����|�!,����@��b3M�{G1|O1�R��R�k�|��&��H�����~7�0�ߖ�����#���'���V��Wy��x:d $�I��f�x�e��۳�j[�s�)MLP�O��*Х�P����	@����Ԋ��D���YDHF��J���e���}�y�hj<�g\)���jx�ڂBgC�x�r�:��7O���I�?:��W����A��ۋ̻uH�W��W� ��]�����yy#V^����*8]�Ƅ+�E�|�}/�a��xj�����N,s'�-����@E��}Z�J S���t�V-�?I{���gnY\j�����?IAh#��'�9�l"A�h<O���$)G#�j<���S�l)OJ�(�Ua�H  ��IDAT�U�7�@js�=}��N�~O��R�5i�wP T�S��=ͽs�y���`��+�#�o��
@%*�yL����T��*T����H�|ޛ�@���T�׳��ق^<�%���	�/�A���q�����E�
>�>�5��� ���.�?��P�}1
B�h�U�cdQ�|�_�|��x���H<�#2�у�`O80g�d�#�١��
@�k�p��O���?��_�a�ހ��>���#P�ӯ�����%*.���P�#���	�0%\��Q-�q{0���nc����ka^�6垰#P����"��c����B��(�7��w�aFv0�fz�Ke��N3 4@˿ʒ�T�NU��,�I�Z���Y��U����@t%����I�"�����7oh ����W��ă��}C�a��D���j�	K1���V�
�M�XU��%!X�!�{�\����<W���:|'��S?�^���D���mˡ�0h
Ӿ&0�nk�V���
@�B� �N��!|���hD �j	@�Q
@�eТ�0�iN ��3z�r��.���QH>��k���h�l�B�+���*@�٪iX(N	����Dz+ *^P	�]Y��Q	�U}J��>�[��.�3HI=U������)��S�_�V��I[��m��-ag��[�~GF$륧�Px��'ːy��*B��lD����/��*����u�8
z]�`h����#(8q		�;!�/Bxt򊫰�7�'�w���1q�B�;� :�����1s0|��rX���`����O�Z�I@�䌙s��bM"�<b1d�|2�B�!k]|V�b��8L��)�Fa��~<�����#a��qX�d.��9b��;���d�91c�L,p[�Np�p���*D� 4�������ή��Љe���#��!�&c�lG��L��2�p��Z��N^X��f����bat��%�爹�Wb�W0�S3����).��s�p���N��1�v���o���Z�\&`m!�, �����Hܟ�߃ ���;|/�j��b�+�
���OH��gG�m�T��P5��`5
nѩj�lIUPP��@��xaa�'�* �G	�� U!��K%|��1-��<�� D׏�˯]F������̽�㮕c4��ᷫ1�v�J��*$w��
��T��׫�F�^�C���Qv}+6ު���q�����~� >��W?|�>z����-�B=���|��@z�v �>�3PH�J;���9ЬF MW���hS�|
�
��CgSi�}PBn%L�ג�Ŵ�n�h*��$�M��Y>m�pY��d��#i���ܝ狐�{�&T�.@�B�tbvF#���Q�ec����HoHF��Td�O#�g��D����$!�dr�� �h��:�8�iT�c�H��[P�9 �|^A��@�%K���H<��J`S~3Q���ºh6���-��:��o��z��V�#�0�<#xL$����(����U���iYK15�	S��r�br�3��PB-r��g,(q��2W,X�签X�+�/�t�����(yu'¯Vb!����;�Ѕe��u�$��p2l����
�%lHm	���G(�`���T%��j���K�gT�q�	��R���gU ��e-e�ms�g�<y��	�����z��BX)��jYW�wR2B���ir&K� ���'��O�M�F �|F5N�
2i��G�Ư.�bY
|vhL�A�T_��&�q�`�Q��)0�jL�Ԃe��:������Z)zݩF��U�r�L���{<EHdD#[Bje����x�F�i)� ���|!M���tW:ݑ�|d��F =��������4���^�eYѝ׃ Џu2�@?�J1���_/��[�zy2�ף��èy�4����9�mo����'���q�~p�N���s���ӎb�kǰ筳���5����.vr����H��ᗷ���&,�P��g�0�ߍ�|��\�G�K���ru%\vay��@$��B�O����@�@��3)^K��R�KB��C�H �-����Q������ ����IO!T �j
�O!�R��ܯ�����,
B���=��D�o��%�׆��p�F=sJ�m�PN�?y� ����H�d��v��g��m�.jۘ&��6|�Z���WI�~GѱgՁ�{�#�ϊ�@��Ϧ�f *�*�4D�<�`���E`�7��%�����V���6�jKl��v"	�h�/���h�7m�vT����Bh�� J��P	+��WbX^0��{_����;�����u��^��l�-i��%�\M�Ƅs�-�4�o�Ĺ�������/����
y'�1)������@���?��W�cJIz�C�M!0��=�0�c§�`�l��z��F�f?Xm�ݖ �s��M��U���wN�{�����?�Ǟ�1=- =�<Й �is(�7���d�m�r?ؔ��U�/����~A��i��g��8s9B�a���}G�����O���/���!L�wCO����.��0�Y�G���̪p,� �UF¥ ��c��� �{sQt��+�5N	K0-`*���.�=�c5�;�N���v�fE�R}��U϶��J]�6u���C��t���>۠����y� ��HǤ,z[����
@�'ڢ�ҡ�@��5�G�͍�XLpwZ�e�zmP�����ϧ�Bp@�	y��<d�!�m1��H�	u�
n�F��ܕ�Հ�h��ދ�~�RT�]pm�=��T� 4B�Hў�)!���h7�Ɩ�;���w��M(>Q��#�� H�-V��?���	X�%��AXS�����4�/Y�_~��O)�އ�ȉS�ڰ��U��Qe��t�j4X�n�ѩ�`t�1�݇�W�qp[�Ș,\�a#	��R)�\���K��P���MX��Q���I�>i1�=Ñ���p_,_�nԼYS1i�H�:Ç�0j��ј9k2\ݗb��+\V��s�����c��$L�3�p\��Z��nK�t�3\\�c���b��3�`��i;y&��P�m7��cҬ�4r
��A�t�¥�;q)����Q�a�t',_�P,[郀X��9�����������0����QG�7��_Bk�6�d4Vx�����������j\̀]��� ���$v;�w��E�sݶ0xm	�'���x6PW tm��P���A�6BnU,��C����eX�L ]�z@[דߝ�� �o�S�3W��s��"})֝(�t���� D�nU<+1�Z].ǐ�v���Ә��Z%��a�[GQs��׶���n4�h:��%����o}�O>y�� ��
���!��M ��}|w޾�W��t>����*P�8�R��+ �l��+�L M �<�"m�gS�¨��+���{@��kʵ�T][���P��p�I�d�L���{�&h��>s�iR�������QwI^�9!30~�(Y�}�wC�Yv�1�z���{ͱǀ=0li?�v�	+��{��?ʫsW"�b�����F��r��/E�4�uϺ��C)a���D �F:7K|�.�Py�6[�<�2Գ@��f0�-)L�t�� ��)��F�M$���	�'�Ac݅�%�`9#�<U��=D���QX�!Nū1���,g��v��\WB��S
�1�x��s���@�Y��\�,Ǣ�5p��cC��;"�߱蕍�zu"n�`�q��\�a�z��|�l���`<�hX�O�9!P��v�ՏӒ`jB�̘jr,&\
�J_QO�c������~�I�\1�>��Ih{0�P����#�4�Db��I:�SBXe�w,Y�R+ ����Fm�+ U���B>D%ݔ�)^j�}�z'	w4den�������
�j�t����s�v�}��+yH^2ҭ�էd�T)�@�5�����I�фedJ�#)r�E�m*]�g����S)\g�R��X�E��R:�n���z�Z7d���$%9�e }�jKu�=�>��,�p��D�n���{kb�nC���(z����7Ob�@�}��ŁG'p����_�G���h��G����q��Q��
^����>�#���=\��	.|���}E��"��a�\ہEg+1�d����@>'�	�=	�=(���@���6�I�uK�ȧ^��]�n��@�J�P��:�-� *����5�@�?�)�
�"�ç��T��{X��I9�P,I;��SI� �B��Ч!���i�����T#�-tj�Y�d]Q�垙&e��x��{(}mۨ�ISǴV}(5}6�J�r��-I��>w>�/�-j�|o��'�@��xj�������@�f�!��|��go!4�&�
|��>/q�% m��й?mB	�!Jm�v�!Щ%���aT �#!���pX4�Â@1� z�������o4�?���=�1���Mx�" Z�F կ���0X�yb��&�~��o�������ߡ��>�'f&b�������~ƃ��B��Ә\�>���hH�4��-0�H�`�:�_�M����¨?�?��M�\�sC��#�?�˟����|���/afj z&x�KY �6��v}0l+Щxl�}a[�N�L���
��_��R�� ������3�J��?J>��+�~�}�q�踌�y�|XF/�u�#�F*˂�XwB�S�֭�C�A�����D�"$����՘~��g� �v폞�{�ۜ����#ma1�,t�I7t4�C�vh��Qk�שU������]k�n�
����o@��Z��3n�A��`���k�� ���At}<7F`�0xl���p��@�p��zI譀�fP��Dھ� %�B�)h�wg�&ܖ������ �����)��eSY�9���0	#%���&������݄U�H��Pp�e'�Qqb���y�
��
�}� �Ќ���<V��3�C��x�C Aȫ8��&�����1�z�Ʒ?Ȥu��_~V��O ����GN�bs-�k�!>������0q�L�����LO�Y����̹���1z�R���qӖc��՘1�#'��8_̘�Ʉ��c�c���W����+��"x�|�z��q̞��S&`�=|0�뉱c�`��	��p^��]�a΢�>w*�̞��f`���J�-�ϵ���F`A�? �OA�����Y�����R�5j���g��c����3p*ԁ��	�h��ރGc�0�ғ1{�+̞ �!=�kk�62�Q{�K�E�d����/��`>W�������PA{7��)!��O��㺄J�)?	������F��P-�n�:�2�����4,�+K ���	�."�a^���-S �^��"��"��._��ek)O�)��W�'!v"��f��k����N��t�
���c֝G�~���<	���>F�b�X�14���Ț{��/oGՃ��S��w���4�~p7?��W�x�ǟ=��q��C<��|�e<y��y�(5�Gp�����%{�ې��se�h>�O�p�|��f@3|�A��T*�P�H@� t�>��)Щ�*a��§H��
p��TB��z꺲�D�L���+�p* *�Y�z,�Z�Bi���ce�+f�O���0`q/t�a�1�����^���60�fC;�b������Q2����Ժ~�V���
�M�A��Kzc��,MX�~-¶�򃓦<����r�|x�+� ,
�C�Inw�G'�E�Ԫ9���+X��2��LX��z!��OJE��}�t���	�2<x$T&J�b�1<.��m��g?��k�8��s�cN�;fd/'p�b2�'�ќ\������^��yΘ�����+�����~Xޙ/k�~��4|���
�Y��G{�#ǜ-��Y/u��a�?
sJ�O�D �9Op/�@��}2@�!1���
L<e]���q�x(�J�g�d���4�D�F%P�j]�z�8��N;"�!!O T�ӔF��ު�\�iw��k�k��P���"�V	ﵹ\����Q��<�hp�WRM�N#W��)|6Җ�s[B�H@A�e1�u�Q�1�Ej]�w�@֥�,`*���oU�%�b�Ckw�H`7��-�T�̧�$.��A[ �P�{&��& �%ܖuB�4���屧	�	4�	�- �s}@��������x��nTa������w��Q�=h��W����Gq��1x� ��A�Z�\���aUwy�_���j�^ۇ�S�Q{bv�݁]gkQ{nj/ԡ��a�yr�>��?�������wn"��q^��ӅL9S�gX�|�e{_�EwB�L��h��Y�Ƴ��x�o)0(���*�<�%m���)��RS��sІ����3��%��,xj�x��s(���!4�)t6�S��|�Y�0Ֆ��j��jҞ��h=�ʓ٘� ��Oh�Pܖ@��������)xv�:a��?�_޵V����N�|��H5֭�ziGX�i��@�?_$����>� �����x:[P�vjU��gK �n������.\h���N��F�����}ah����цj[���F � �P�mw�PiZ����	���%a�?��{�����������EBw{0���&��۳p��'���� �u
���?���ޘ����E_��K���T\=�I��OT�� j�%P�p�?	�F\�Ѱ4�]��~0��Q�h���z?�3B�����w�aaF$�E�bXVV)��u�TH�-��q�`���6y)^JY���h��
�W���ܬ\�豚G�׿~�G_}�snшMF���z�0��:���`� ���p����]X]��@�m�Gơ�7�!�@A�i�S�*k%Av>����`���b�/郮s{�Ӕ��mG�Lc�L{ڠ��!Z���%B�����VP�:�F�|� T�ۮ�j���#z`���h �g�D?���(�C��L��j����X�1�5P\* Og�fT\�T;�S ���x@%W#r��s�\�/� ��w�
P �,�2m˸c��m�'J�_m�v+��PQyI�Ye��S�X~���ʓ���){2���d�NT(/hl}:B��jhG�%#lg�KB�kFt��EO����6�؄��[����}G���w�Ç_|��?�w_W_y5��U�U��b��+������#c&,Ƅ�Θ0��F-�8.�O_N u��1K0|�+�O�4�m��0}:m��K�p�2�\��̓��9X���χ+�u���b�uw�*W'̙<��M��#0i�Hjf8L�b�X���	����3��X�t��\OO�\��^����$�.����0p�h���gq���43�-U�}.q���I0v�#&Ns��"6�&���Y1c�R���������`*l������zN��ÿt���L_°���>!|�և!zw��P9[�;����!j�@q�P�;��+��n&<n�Ǫ��X�9P>$ ��d!��]�<����@��v09GJUnXuJð�4�e�X���]����� в�tu#��4��W����z��)݂�s���|�2�T��}��	��Q�+0�i	R�/�cΙx\ހ�;������a{�n|�2�� �}��}�*^��.^{G��.��
^{�e<|�.��*�|�w_EÙ��ۑ���Y(8��4���̥���éjP�8�㈊%�E7$#�>����U�Bw:	Ea�	�ܖt�/?	όjHR?�̡#뚼d�UB�3JDT}2_�4��OGܾt~\x���og&�(�Г��?���x�xCS�{*E��QB����q�QpMu�d�	�5��'��v�	̇����r �r��F[���N�>����E��v��(Y�oOuF�q�g�-���A��V�jk�a9�6#�a7��gv�0��p��P6&E��Qu��g�� N��#��z��h������@>����5W�xFY��k	��W���74�9*/�H����C����i3�
�� �oOt��Aʑl'�]��d��(%��\������rO8{`q�r��v�\j�Ӂ0:+���pN�tQ���)"6�3rW`v�*8���/�+���
o�T����X��k�	����e�~���7a!���4~��G`��d�>��^'2�C��4d-i�ڞ͆�Ҋ*�I��d�91�w2Uy�g���G�4�Ұ�%�I�L���' ��Ɇ΁�싇.C�'&G	W\J���bљ��v카"lZ:-N�����k��P֗	�$i�ʔ,���<^Fݵ�slC �`yM�j<��4,�	��[	�r�=��V�њ���|:Z"�	ޏxj��-���ԜH�1-���ҘF�����zު@��kГ�l�:��zF�3�Bd�3��އ�&e$a����r��8��O�� ��h�m�'�O������`v>��`,]̄� ��\X\�A'�U/����x!���`��D�߉�{{P��~l�������Pw� �w����C;��~#6�݌=��Pj/]8�[����?|�/~�~��{�o���S��=����a߿�6�fO6�#�߃������I4�~�OΣ����oq�˻�~�
��b8���-��(PS��|��2�ʕ�\͇�X���KYлD�:�'D&��@h�Ӿ�M���)o�s��ߵ��j����ұ��%>�����j��t\����u�i�����6W>�m�.��<)��r�=߿�|��i ��g@�#w$��1��K�S8���;�w���O�k- ��vSI�*C�?�$M�)3��"�]P��kכ�5��j�0����H�Q��}�&4�n싩D���6e�Y��D;�fS=�w) ��'L�(�8#X�%H6W;����V��ю چ��}�7AP�E/6Dp�Y�����}^{B�b](^�،@��Qjࡗ��Ҟ@�jT��Ԯ@�����Ξ`t�AǺ0���.�a\	��u_��On@�����
�1(���ס��0����X5nG��Nm ���æd�oO��o㻿~���O�+�?��Ѿ��o���L��y�O�w����eA0�	�ц �Pf�a*��aDC�dS0,�n�%�4D�7����N\۰E�����'�@T��`��K������0�4P���FG�^�j��F��h��6�K�.})tӝa��6�a�=��X@ ���#��k�'����8|���b��(�~>�0.u-�=��b�8VD"�p9��� rg&R
���I;ӑY����5�9��R,�5��L��1�jz-�.s��v:�s�=:M��Q�`��m��������Z�}�vh۞i:�zA۶m�6\oC0mK�!��o� TG��j�,�Xa��du��������*7�T|6F�C �:X��T�IX$�j<��4Pə �\���\��<G�w��h�\�`Cn�� �����=���Q�ܗ���H!��NWN��a�-�tD ���rSK[jG,����L%��T��t%
��"�^3KƁ���VK�u����5�;���̣EY�޳���.:�5��(Y_�� ,&��x�@db<��lƍ{��叿�	���8	�GN`ߙ���݇��tL�K;l�+f-XEu���s�w�T�;O��5��-���;�Ƭ�K�d�
�,]�y��p]�5���q�#�L���c�c��)X��gD�!>��������B��1z��cǏ��3�p69`6������E���m������p�Z�G��8k6���ai�&;�m�/�{��a�r�t �-Y���c�L'L�vdB
+�!��A�	X��π�Ⱦ0�3���Zul�ux�2�7��>O���D�ٓ��3ň=��k�}>��Kxm�d��-K���-��5O%�
����<f��(�?<k��99Ǌ�w�1��Wմߋ	��AX��%I+�8��p� �0\/B(Eyu���K��t�Vi<�2-K�7|�}�W䅘� dW���x����(<�	1��g�0��4��˴�E�z�0z����c��\�&HM:��Y'��X<N�#��vl}xG�9�����o	��>�~O�y�'_>ģ���ỷ�������/��7n��[���� ���e���@Ѿlh4� ���#ҿRF��J`� �7�PBp$tH�M�NAG(��-��M%���#��c�y�v�%6S4 J���~��C9H>����T$��@B��q<6�D>6����*����'fMF/�ΰc���2�]F5j���GX��H���eWtm�.#:�n��s�2��Gأ��.�=�+��펾��]�{�=z��幖�f
�a&�b +�@���nV&� j{4�s����y<[^�;�u��c�I�n!>�;	�;c�*�����B�p��-I�	��GT�C8[����(��b�#K�L:���"�|��{j� ?�X�k|�Z�
�
ݱ8��s�c�@(�y�n�O��M�X���t�g�&�,#��Ñ�Y��9�P�O�-]�Ee+��r��{a�?������w��R!V�υǥ|�_)¼��w(�bѝFW�]htv9��N'3`%��Gr��a@Xԣt��K���	'aN��gG�h�u��ׁ��	���J1l.��$�y\��V'��ٰ>F�<�#����S��`M�!(Z�"�4-(c�f{u�}lK#V<�25�&$�G�7V���WW��N}�e�����	�
0K>�>I�j�O1vi���` ��S}*� ��Ic[�P`D�����W
��Z1z�*G�e��\ C�mp:	���gh�����T�v��q����q��j8J-���	�r{��Uxn
L.���|",�'���������r����j�/f�+�g0����x)޷�wo;J���G����{;�D��E-��X-��=��W����+���e���[��ˏ����͏��;��G��'￁�� �|�1���w>�>����y7�_���p��!�:��O��V�[���f���P��A$߭��M���$�/����Btb�Y^og�/K��L5#�޿T�S��� ��K�!���Ц�'Oes����b �|�l��m�;\�y�4�q��5�Q���uJs���=hAP`Q;߭�B���>$����|�4��Be[+-|j�L���h�鍚��������& ����w�,	��u�+���ܯ� 4:��ͤy���	\6�L��#`J Hl��S�C2�'���s_$��_�$�5� �����/Շ���0�j屄Η�Z����um �P��:�T;�c;.uw�|C ����k�J�M��#�e��G߸j��^;�`�+
�uQ0�ׄ���ͤ�f�#f"�\��?��߿�G4���_!��`Z�7�߹Ĵ����?ǞW�avA��z�WY:��%��j},	<UA0'���'�VJ�M?�b��|���jo��[ ����p�0K�+�������X��Ѯ��kg�'�m3��.�3�a��
�ū`��
zqN0�p�i�#V΄��L��$��'�) ��W��ǯq���y�>�uޥ.��.R/�ĔL/�Z瀕�vzR�����fl�Y��Wv�6-E��l%�iw���đ�0�<F���.	�=a?�+:��N3��|�����U+����m�T�mu!�@۵!xB�@۵'�>۶{����Fm�c�}�1� :}�lt��Nð�*�j�9��B��p��	�u��X�ɹ�Y�T Z��U�5��^�	�k�.�)��� (��	�)'�L�S"�$2M"Դ��2�I:m�<�E�F�v[b�s��u]����<����4$�NAھ,ds_��<��F�k2g"�@&��U#jK2z����z�7��<�WQ���P,�Z���]��Y烔�,�8��W���W?x/��v=�Ԣ
xGc��5�=�ash�-��b'?,Z⋱���qX����289����0a��p]���X�Z�Ύ�X����27,[��}��X0g.&��Y�'��i)�����I[n��Κ��3�b���5jƍ��S'`��ϛ�4� :e�4L�7��̅�w��B��������]0~�L5�'� t.�"��X꺖��"�5X����J��d!(2�e�Q�a�2��d�*�[:�G�S �����;�E�Vhe�]������O��.e�7@SԘ*2��7T�S��O��۲|@	�^�้�1@y0��[" Zx��[�V��(~��X� �d8&.�s�*���R ��T�O��ju�@WU���?�|�=
$���H/�±s����;�Pyj�.l���b������eXy�
�o��*j��J,�R�e�K��j|��G�MH���^?��^��o���O��oo������x��kx�Gx��W���W�������q��۸��<��>�_ŭG��pn
w@Ulz��3�j%�P��%�
����\��ZRLC*��T�{�O�Lo'�S$�-�/jJΗ��F��2��'z�F�y]`9�ƃu�Hm��uC����k�a�N-{6�[���)l������{ä����7�qg}�v5�ywcX�2�m_Kt�G0d���l�k�=���;j�`?�6�Q�A�,0j���1?b>��h��OG�<5�n�^�.~��`F�"��Q1��Q*4��(�Bc��7������I�dz��ٲ��8H8H�����Y%`_0�JO8��Ҽ�X��E�<6�s��0���({dB�<07s�a�) �Fv����9+0#o%fFg�$���C1� �X͏d�t�����������Awj�}�J�G3�g`PCz�A�#��Ip��g�eI�4>L���{��'R*�;�ڋq��th܉&��HH�3��eA��Qu�]*Bw���ɨ�Gi0��D^'���%���|,	��4�L	��]S.H��F� �\H�<���0^#^[�S��ks0N�Ϙ�J(��8�A-�Ηh��� �!e�J~���
�
����n��S %HNgB#߂ƾݥh��R��w*������F�x���c�M�$x�N&L�~	�#�ڎ�lG�[���Gc�1�w����z��.���B��iF�4i�H<�2�!��2��0�B>\�W �A-25���!l��������~��N���;������w�۟��/ɼx2��o4W�������_=�f��M�@�Q��x^���s�Q�Jn���jGƫ{�G]~�
WJ0�|!�Y�y1�������oFI��@���/!�� ��O��J���i�6��� }
���j�������\ͯ/j��-��o�wB���wF�� ��N5��@�O��SS��� �ڹ-�Jޝ���i,��~6P�O��Z�͖$ ��Q��=|�Z*$X����7�=T�JT���xB5�:�v�7���L+NeS�T�h�P�6���P�!^���i`3�y�!l6�D���{w�S�H�$K�K;��j�Z�$�6J��W�`W�%�o�7�<����fʀ>o���hX��	�M��������u^�����h\qwww�	�����$!�O���PJK��T��Q����^sr ���~~�~����f��3gΙ�{�묵׎F?���~|>��F��n���ߪl��=�w��o?����=�]?�YA�X�B ����?~�{??Ğ�2;c�\1�,�h0����T�K?B��X�$V��3h��q�-�\Ӊ0���M('���s?�w��o_Æ?�	5ǨLg��3� �Z)���b��Y���n�f�N8و6��a�"��x�[i��ǉ7n���?����O��sx��p��(}�	���1��� 煰���K����@FC1J/�F鹝Ȫ݌�}�(oaH�X�l;�&��Ř�3��b��q��Q�Z1���G��}��O�>�j� ��'��m؉�k�.ûa��b�ـ)6�0�f&���D�O�gy�3T����Ax�I�a�3<����Eފwӽ"� ��O�����*^�m����~o� ;�?H �ag2K���g7��L1BwE"�&����w��ِC0�Gҕ�h
��h�&��=��Ժ4��W ��"�go��ڴC'�L���3"����{wg8���'( ��
CBR*Rҳ����=Gjp��p������=�;���"l��V<�3�b�����gԄ>vb��Q���/X���V`Պ�pqpG�!����pvp���<]��� ?x���r�9�.X�y3y������D8�G[k�Z[`���X�|	�-Y�%&�h�\B�|,[f��X�n)�X����c	�t�&3X:���Ǔ �Є8x�����+7X`�ҕ��t����G 6�xm�}��a��7띑�[��G� $=|�0�b%�͙ ��ݡ��:���ޠ#�{�a��z�zBC+��qb3r/+�r�e�������i�
?x( �C Bs�ۓ���0�n�w^\r�a�쌍����p��f§��� h���.%�3 ԣ��ވc{H/��Y����[gQ�jv�Q��{�P�n�|Ѐ�Q��1r9�u�!�#��^-��k������~*_>�wkP�z��ք�4�ԫM8��	\z���w7߽�[�\��w��曗��J��>��x/�}	G/W��0�p�۔�?P�@h�7T��'��k��X�k6�V� ��TD�RQ�@���d0pa��|v\َ��t�Z�8MàŽћ��wvW��C��6��Q qa����0#t��>����,.�ІN-%��?�����k)2꣋n�>ûb��^4��9�FH'������1lF?���ݦvƠE0�f:6Dn@ ;�ԣ�� �'��̵�$�YRwsy�c��j�g�ߡ�Ӫ!4��/`�Z
�r_�|*a�
��:��L��m!���)�V�ABC:��ʺx�U��4���q9�y( j�G"7��k���8����{�"��|�n�p��tG�)A4M@�KB3�o�I�e�b�fk,�6W��,��Z60S��rl��M{C�T���T���A��|i�.�c1asF]<&��a4�o(A���4��*Ob��&F�5�&h5�A��f]�h�u�k���@��Y�C��r8�lԵB��Y��7K0����R��/�T4�P<�|.���P���c1k�`L��F#Z�8����K(�,�WG���J�!nO����X,�&n;��6§zRy�r*�4��x�c��b�7�2�[zaT�)���݈�u����2�r?k�Y�BH4<+�>OƪJ����v�<��F?Դw*1��J�\�����8����!w���z�r,�ʸP�8Q��J�$�%�M�g]ue<_ލ�k���Өx�$����k��>{N��Wn�#�������;��������w���~��7|��'���ԞkĞ�Pq��V���k�w��^��+�`z�O�`�����2�R�\�FOJ��~!WI:��|�c�l)	�(�7j�j��>�� [�� ��п���d?��S�gH ���zy��� �ܷʽ��PU�-�=��5�K��?hK����^ZHK`Q ���G%,���+�I凜)�X*���k��J��Zܦ���W쫤���f+)��}��}�Fm�?J�G�T��	��@Um렄��!,	���n@���R���{Jm�v��N������U>hG	��g���P��;ap�3v�{���~���x��q��7p샻9W���.��;�0v_�~�-�%{`���x���������퟿�=|��Ob^�+f��`��S<�������_a��X�G Mv¸mA����z������9$�i{��k���`r�'FG8���)t�V����o@��C���)������޽	k{\�9���8��}
\ѕ6M�t;��pD�T{t�������cfb(�d&��b+*�\Í�����p����Ż��p�+�~��~Xd��.+��bz��B�ih�t &��Sy$���V���BN
⩘�x�Vي}P�>��-�4r�`��,����Q��cĆ��f.�A�B{�6:�{<�� TO_:�\'��i��ӆ�?3�eX�S�fc}�-����s{�3Ԏ�)�'�:���l�W<�-eC �)�y�u�g�P\G�T�6{B�΍ǉm�D��-�?���d�U2=G����1����3�x$MK��$CÊ�N�L��VJQ��,$դ#�
��CԁD��J�=�x4���%��N���0��M���5��⑐�H�􃻗'�����`�x���;�ˡ�ONC�8y�"^|�^����8v�:�2�`��LW2a�2,\i�1 Q@��Sc訙�0e&Q��.pu���u�XCг4�K�p�����|�����%������=������=�������p���j��
��r��XF�\<.Ι��sf`)�s��%Xc�+��V,��e`�z)�Y������1��JC@\4�<\�d��ή0��Ǭ��1r�L��.�!�}�(��WB�x�`��e6W�ڄO����~h��æPk���B��D��S"C[�@ś٬�@]+|x��(P�m�ܬc�(:��	*&`�І/��+ۦe
�^�ԕ �Wާ�%^�NO8@�J<]�	�n[<�S���?��F���chS���m�����/N���Wq��S���	���;�=������}(y� ʸ���C��w�_���+;Pqe��Vb���<�{ϳ��6e]��_���K{p�l%�߇�k�8����;��ڧw��{�YW�-��7� ��D(�� ��Ց��'*cB��%���œS����%�S���#�Q*F�&M~{0�SQzy��ه�]�0q�����h�&����й}1j�`�"tJ�젉�L_t��޺����F�iĎ�3;Ec.���4�����Bp���릥߰�6�2Ā1ѩ1~�L1�q�G`���i2�V��v��	�����qlB(�#I��u���	*^d�^���T �.�%^���J"�V��4�6��������4�أ���яDh���6&¦��%]��"O>�+y����*e#���-l�~p���e�+֧9bM�V�ڪBs	�&�6X�a�9V�%!�
�sl����f�ֳq�e�+�|@T���x/���R\.��bVK��LL>��������F�4�A�K�L	=kT͍�$�`����H�G�[c�F�(Ĉ˹FpB8r>#/�a̵�!��"��z}�ܫ��0��"xa�Ļ;1�V	z�NGB�!�B����M�GCU P�F���*%�N�v:FÒƨ�b�'Ø�ҕ�&�:4�o&_+��q	!�A���>��:Y &<�P[�ӐF�Օ��K�f�;��璕0[�1|},��$V�=�E��q�����v�1��Iƀ�يG�+�Ԉ�ip�b�����8
�ʸP�T��3��|:!6����ݙ]/���{���r�gWp���������!T?����������R��/�S�I����ן�?�^����S�S��8Г?���Y����������M��N0n܋��]�q�0v�R��׎"��^؞)�򓹘u>�/�`��l��zʼ��e>�<%ɕ>�gK�T R��Vk����>Ej�]k=@��Yj�k.��N�����Tm'h��
\��jS� ��!%�i�N�g �Z-!T�>@�#���bG�í����T~�Wb�V��^�|O%����������>�)��I���&P����l)��k��bߦ� �$!���A�!
�^ن�����mm���^$���`S���*2	�J�� ����f=�ϗۚ��ܯ=!T��^o<���+=����4��f9!������|�>>��<R<�����VY�Y�!����a���~��W�k_}@����ǿ}����c���+��(����Pq�$���/�	��=�<ӜP��s�ز@��O���]����D�Bw��l���R֔�?����>G���O5�Z��N+��>⳿*�??��+4�vV��a�k0$�C�]1|�/?�+"̡��nˠ�׎�]�/�o�.��&>Pư������w/��k���M\�{	��X�k�~���p�0t���^.���m6t֏ĴSؔȲ}a��ϢP�W�#�*ѕ|�JE��d�UƓYf�`y�j,
Y�Y�s1�~*�ZM���	�Q�1r�h��B��9�*j�	}�X����ճQu� �NnźpsL����I���2�3� *੖�v�l�>�* �\�'���)a��"�z:��C�S�	�zW�#�D2/+ *P�m@�Ǔ\��]א���xe,��f��|�hR범R��Oȉ?B��vu���^Q��B�F#�d��b��
t��Cg����-r��"%#�Edd$�#�B0$�8��́0��G{'�!99�����W������|�g�!-�~!�H����$�Z�~��a��)����;�K;��8������ݸ��noogl+.Ə���<#� ��d�a�!\�t�ɉpr������7b��)6���|�Z�-_��bь��3e2�͝�%&s�r�	V�[�U�˱l�R��"�Z2�V-�'KxD�ß@����$%������-��
���㘮�T�w�D\~�B}����̗b0��nCzC�+�X�����&�ɵ�nq�u M�u��*@%�!T��@�*|�ӗ � �9F~�(8Y��r�TYbvH(n�6�:���a���|o�E_�w3�������� �R��|7Ĕ k[,N_n@���e��Kx|y'!t?�>>��oVaǽ���J
n�!��d^߂l�Y,shP��G�l�ނ�s[��B9v�,��E�J5�����|lm*������TƲ{������ۍx��u���u�^�|~�y�����%!�h���MJI��׊g���/�J�O�� e�k�h*��T *�T��e(����p�������1�y6��s�zO�ǰ��1rN?%�v��~�?�7z�νa�UZ��:F�FJϘ�h$ҁ���Q��HK_�5�m@Pm�l�RK���j]��d�ZMt�#Ԋ�#v�]5a�K=vƠ��1� <f���;���xv�c���D��X�f�'D��sfߌ�C���������'Y��R�
I�h���S�
:e��R��i)*�0�%�
@��* �z"	��ī��h?�l@=�����n��pg#�(�C@y�+y���+�_I(�w�#���rBiQ�a������a�KSm�X 4G��X"ʕq�X�c�UyN0%�n��ߒ�Ѳ� ���lضU�p�����\^/�ew�+�fcH��Doɐx8�G M��S}$��E���p%ɆfMtj��{0��0�J&�*V��tJ�y	X4`���${R{5ġ[]<�7$��Q�Q��J�1��0��g{zcz���]5"�vf��1e@CӐFkg��iHk#7��l�1I�_�Fi��Y�y5Ƅ=���ӣѪ���Jx���
t6K�O�"F8���*���k@�Z��rg�!i�� hw=K =�c10&L�<���,�#4v��܅Fow��@hOhϳ)��t�;�J���g�$�
̊$�W�|��{]���~2��f��Z	|n�F�k5�~p��^Bեz�?W�s�����o�e��M��P���������Z�^R�����P)��7٧y]���z��°�o���?��^}��]����
��܍ݷ��?o@�Y׋۰�R1f^��IjEI��^6����0$t+�:J�lH�f�Ԡ$є�$�!�=�zʺ�T%�o���y���:�%���c`$T���R�\r���g�} U����x���^��ZzJ�xO��C/����O TQ0*�>�.O�n.u��O����*I��N�ɱ�㨀�)�{+`��֑mP�8�����%�M���J���M�WM��B|?��*��I��h$TRZ,��2��d�� pr]�e�ҟu�vu�V#�C�����XB��C�d]�V@4��4��؁wJ�#}#��AI$�鏶����%!�����6{|X��m5!�Z��� J�������x@���{�щ�A���B��~�[���B�QW�o^Ɨ���~Ï��O�0���G�^=����j�gIv߻���~�O�	�I	���p��:Z��F"��:`f�-��9�o�+����C�z�11�	�s�1�,��C0��3��tK�à8{�J�B�����o���Y�o�D�u�0�z)���"���G������5+#�W���"�.���2����Eh�9�AX����:���W�����z��o�����{���[����㣟��O^��3���C�L�h�E�}�桳�t���E|�:�� 8���o4�3�:����I��$�쉀[����2~/�����<�a����0	c�Oƈ%�h�JI"M§HC�"xjSZ\ �lP-���7Ң������c�ڹ�<�)2�:��1��W'=	�-#x6�A�q�ʃ`/�I���6�TKY���[��J�VPe]��P]x���td],A��2���GT]*m���=|��Q���9����td�(@�)��,S�ژ��{Uq��dZ��F0�S���`����i���)rV�����A�9�?�,�#�0qIq�GxX�}isy�!�'a���s񆓅=!o=6�1��zsXn����+�SQ[ӈ7�z���~�_����^¹��{�o~GnA9��\�ի7`ݚ�p�sB�o <���p��k�u��d+�������оC��·/�cGy%�ܾ�=�+�c�64=��#5(�ی��0x�;bӪ�X�p1�̜����i�`��ј=c/��5�c��X�q��[�9��bΊyXh�k6�+��+�Q��r��?�9�����!A����Gl8,ݱ��36�`����9�t��BG�a1� ��`�x@��p$MД�9{[�P�PޔWu(<�6C(AS�x+�NPʭR���^J�v+��I8u)�7�ͧ����VD�=^���h���=?HP�]����u)&\{��X�NE.�wg�\J]��D�<�3md�B$�E~E2.H�R�ds��"�x��/���v	�_چ�ۥȽ���K9H]�A��L$�xLhH@jC���ϕa�٭�v��'���X>
�~��S���<��m�rT��D��*��<��_�˟��{�s(��)�9!!�� P�g�c UyAE����SA�Z� U<��"����*����)�T{?YL���K#d�㫎E4�/jr���=�w"�<�fcؼ�9�'&-���bЄ�3�3�0V�Ӱ�.�u�'��'E�4Є�Q�u�u�����z�>��c#h�,	�"m��XzF��N]��"m]eb�N�V��"=�PYR����n;��	��Ѯ���C��c��^;{8�.��)+&b���z<�;.�e�"v� ��׿��a~��b	��
�JG���S�<>@%�V�RHU{?%��z�����^%���j�T��W��<Be=���	V���
��m��`'�#����m�%x��䱶�^(g�
GlyR��"u_�2�:`k8ܷ�!��rܰ.��R	�|@.j�-!x.�q�r.��v��fl* �Rlh�`^�
�roسCp9��^'��~v3�h蛝���S�v =��Bo�'��A�!:�d�0h�F�ϹL��Q�q׊1F�m/�N��OC<z�A��8<N{�ǠgC,��d�i���{2����e�7߯�T%�x@ų؅��#���1��L�ze3�}��ICW�3�ٙ`�Y`�F�A�F�AT����$�g���@�h4����<�<�,�]˘Q)��~"Iv�G\�ТC i�5 �!��T��,R$^���ټ��uA�� z>C�G!<��Q. ڋ@Ћpԍ�!�QQPJ �X��*���"du��]��~g�x�6\.���]�|��;��o����Q{�8���~�a'�) ��BaB5'>��V ��Sm�Y	�����y�)G��r�Y��Mȸ[�����r)������Yx.���+a�X���P�;�M{N
�R��Ձ�GJ@M�*�T�ꪦQ��M�IV[5�=K
4��S�R`�q=�]�c���S��/��O���`T���0��O�[K<�"޷-aT���1���H�T{?ա����|y��I)�/��k��l���7Ġ�xY'0)�R�7x�/����iI���%����������/"j�E�Bd��+*�:����>R���F�5� J��B�Á��'�;��wd�F��������_�I�pP��m�z)z��G�sUބL/�/gk<�����5K}����I�T��>;����m��w{��No���52�gv������x��	���S ��@��j8e� �`^��a�x??��K�p�%�zp�'wbY�f��`|���[��S�ڟ�ݟ��_���>��Wo�sw�F�``���a@�+z�;@��["�����|��R��Ϳ���~4' :�Bṃ<����_��W���?��^EPI6�Z,���9`�|�1'�F�T�r�^��?�$+��������-����g#ٛ ~{,νu�� _��)�7�,��7L��c������q�;J	X�i����@>�c�/1���1��ݕp$�|�
��;`m�,Y�Y>�1�kf��#���K���$1���x��g�g3x��6��1�j|vPyAuUN�n�3�bݱ>���	��`��I)Y���b/ JP��&�'�d����:�J�36�.��`*�O����-���$7��f@��mQƀ�����E*��q=��R���c��y"��9\�V��$���3	�«��_������D�h���J;^��#��a��3��hhw%$5�@��@������ށ�	F�O"���i�7[Ev��5������<��[�q����⫸��Gx����ɗ���P#lܱb�)V�X'���	�N�tv�����\���gke����Xo����4 �!���EHP�rrp��I\�p	��;M ��d�e+��dt.L��	#�a��;r(�L��S�aX�t�Z���`ފ���l�Y����`�m��`��D!� ��q�� ���5�.a�����#;�a���a�5�����Ymt۠��A���{��d���U60�ƿ:\	��=� �$#��=E��
�
|* *�>%��}�ǀ�T+ *c@�ϔ��d	��xY��ÿ�p^�47X�:�>[��2h�ȝ���Ů�(����-#�n���V%׿�[�ܝ��x�$���D��0ET��d_��E*�d"	|��Q�|`��^E�����YB�����8�u�g�P|��g��h9?Pɱ2ߎ2v�[OV`��#���e����^��éȩOE��g���K�{&"�V5nS��|�lt���Y~��l�s&I J^/�)a�R��)
;D�0�eʕԆle���;��z=�3�7M��y}0ޤ?���Q��`���0�}vT�:����	]B'��/�:�e��!��P� �=�P.��#`r[K)^Q	a�C�:�Q�P-��d���1e�+M�D��:)�ѓ���L��CӰ-zj���n1m(�-���k�c�ک�f6s���<�Aʤ��YH�IAA<r_�& R�,e�f ;�g(;B��q������XܧeH�xB�}䚈�S$�) *Yy�zʺr=�_hU4���|�U�3��Q�3nO"��R�P���m�WJ��=IIH�NW�E숅i����\����;a]�=Vf8bE�VdQ�ΔV�8be���y�6f;bC�6���q��ް����08�39�>� ���׷`!��a�y���zFWyh�O�]�Y�oڍR�:����R��(�.��ލ	�d�%��a��G�t>O���f+c@eJ�aW1��'c)e\���a},�5�+ :�<�'���E����d�6��G�cI0"���uiD�5DCG<��7$J�������Bg�㾗���j�1F<?��)JB#e�qgɬ+�g(y˝y�yΣo�Q��L���	/�b��%�/��A�17
�9�Ћ��B��N��J��LP1I�.�F��+S�HHo�lo�s���}*�.#��d�=��.��;Wp�J�]=�O~E�N��c2���S\(�����ͤ���M��2���?���^E����vt'v�0-�{9o���}X{���`����~>��tf�o$���>X�,5)�gG���dBe��
>U���Z�g(P�x����x�Z gk� U{:�g�1x\�JH�
<U^Q��dj����O�e����Sçʋ�z�
DUP @�����'�(�����:�Ҷ������?)F��c��T���Y+�a�8"�-��z�,����k���x?	��� �'���?@�;��m�#\'(�# �l/p��GQ�jo<�ǃ����g�d�M���������mk@�V�X-���
|Vz��Ed� ���Z�ܡU�m¨~�'�lsG�\,���c�Q}�4�}�9��������'���׸��������_��_�[<��?ƞ�=���`���^�g̨��ȿQ�����)���_�#�b��%Z��c��F�Za5!ԉ���Nf4���_%�Пx��#���'������q�vX��.+�tl^���Ï��⷟�4����p5�����p�Wp��q���ޣ���w<���l��{|����p��iޘ�~�ZNEĶp��
�<||��5`}�5�l��Q^K��{!�@�m�ad�
�ў����.�g��UɈڛ� h��x�IFؾhx��®��3-�4z5LB��$x��-��yg=�-f`Ԫ�0���<�Oç�Y�)z����2�a'���A��=0b�X���k;�<���P<���B� �x?e�'�<X	�����Ŵ+i�b����MJ�M��,�jo�?IBq�h�&HDqMYJn�? h2�3]�nrhϥ+yLd� hX�b*�@�2�g 4pO!4�'�hR��ç cVMG��}0�d��]�L�;*������A�/��7a^A��DFdB<���Ooyx��ō�hO��u�p�w@fR2*��ą˷������?��k�q�P�6k׬ǒża�ʵ�O��-B��Q�O���'��ly\­��x.�>���E� >6)�I�N�M������j�F�Z�&s�a���X0}fL���#F`ؠ�6t Ǝ��GaҴq�9o*�-�����gc��ل��X�q9��o�k�'B��L��;.�0�r�RWs̶Z�1˧�ߔA�9���v>!��^�_5	U�J�t�(!T~4H=����P%�J�jϧ��l�����ᵛ�nS%!*8[��S�
��D � X	��P8d{�:ݕ �A��� *c@=�z� ���q�{��o$�� gGγ/j�u"y4R/�b˥<^ٌ,*�b.�h0��&��H���K#$���:BܑH%Cj���J�\�gvC.�q3r�yg������(j*����(>Q�Bv�[�� ����ˇq�͋���u�y95�J"��HB��'��F#"��ӭ��	|Fʜ��d���T�F�J.ay}K��S�e�}�P���/���p��:T^��{�3o�Q,�<��9}�g4!�W[hui��5"du	�z��X��iA���N+`*^Q#=�B	�Q}cc�3�@��hI�-��}u�	�F�ԓe���4և�5���R�3�֘��(=�Sz��Q��2d�ڹ{���^����l
���l�Y����f��]�Tܙ���դ"��*�'���hvV�Y[���l�|ʺ:���S^�v+ӯ�WU�r� *�k$�J���R�2N4��.l/��+!�#]���=	��L@*!3�@2�2��#�[㐰#�;����A4���HIB�E"�,\���f��4�g��4�k�\�:�kr�'�%���v��v��a}�;!��)�7ldC����������ap!8���n�Z�S����nuĀA�H�p6��kb��Pz�ģ�1���,�cٗ�*���O��ϩ<��~��q�os��$"p!�ePBVgJ�]h���A<��f��]��:	A,��� ���DH�Ӕ�.G�`XAx�������I�B�R��h����-w�)\؏t%l>K����4�u�F"�0�Z&�\�!�2����,c.��3� <����J\�T��F<����\7�ɲL�BI�Z�	X}��c	��N� ��.�R�C�]������z.�t_>�R�|J^[I�$�������R��!�?5�o��1��O�T�P�N2�ѓ�(޿�Ǫ���e�?��`���u&�O��!<v���d76����+��N�RЁjG U�j<b��-W����{J����*pl-��?��X���S�.P*�G��V�.�=���S�ghk�e�S���T`R9������� T�e�uO�Xu^2�U����I�Ϳh4�3�4(�z�N��K%RC�3� ��!�:
-�k4u	�:G�ɲ�ir?œI�l��σ~h����u���<�xHe\���w���Uj[�E�B;¨H�����{l>C������ R���>�:q�a�S�+:�tA����˅�λ�Ч���]0(��;����Kx��x���կ?�g��G��T�\���}����h���7c|���Y�������7;`p�%�f��3���K��ӧ���Y����k\��m�u���aT\=������g�q�����|�9���{��WPv��(	#�W`��2>���}��_;��	���P�c����Ꮯ��xiŃ*[~������o��������ރW�p� Bs�&��fb��l��G��'W���7���o����H'���a�>>���s.��f���<l H�n�]�-? �|�FT� fmν�ʸĘC�&yJ��m^ؘc��I�2�+�M�(d%��-��٘j?�OC�	=ѱ!�|����g���F{Θ��	�!]0h�p��8E���RrIW���&H�2K��)c>	�;$��
@� *�iWʒ�J�!�# ���S�%ӭ
LU�-��}eh��4%nt}�k��%��� �X��L#G��6�`/�)�F"�h۱.�6^ T~��m"64m���x$�����i��C�bƒ��v�GDR"b��E���#�!ԇ�DBp4��RJ ��������np������`�`WW�yx ���Y��o��o����z_~�->��3nي5�6b��
l�����+֮ZO7��S�-y�J� o_x�\��66���ơ��x��wp���F��� ������L!��gkmww�~�j3�Y�
s��F��ıc1|��Æ��Ic0k�̝?��N�b��5��z�
X�X����a>Hڒ�-U;���@w,q���՘�~F�L@߉�e@��o��6F�a��	2�(�ђ@J¥S��� BhK�#�6{=�q��c?���� /�3t��2����*CԮx�>Ô$D^[x��ޤ,c@%	�?�G�
@�J�����z�z#��	�������&�IkHFαt�i&��e#� �}9Y��	�T��l$Tc��3 ����B��h��C:�S~QI�_FX�F3�Y'���(l,@��R�܉�R�ԗ���N�pM��������Vrks�eg �1�� sT�S��dB�0PU�mK�S��*Il���7T�2�T@G�v�UBvިD�k��z�q6Jf۾S�b��7�3�#`�m�N�m��m$a���ta��C=m�kØp�P��N�J�ᴣ6���`Ե+�������2f(������`Ą�\������~�9�7���Þ�֞]�������E�u5�~	�%|� z����$-�������5a�� �����9�0k%Ӫi��l<f��sI�C��h%&�6Uy��'4�ߝ|��.+�>U ��P�zJ�[vh�g�:�V���J�]�>�
$�H���l�T�%���#�Q��&hV�#~w"ҫ3����؞��LAʎd$�JB2�SWN蕬_�a���H���o���a���/�gz�,�k	�kr\�*�+3�2�k2m��EMs<`��u�T�	���`��hU�	�Rwl�J��Ɔ�@8K�/���V)��b=Aqͥ�0�:�n���}jѧ>� J(<N�<��~'2��t!3=�����t�>��>l��+eoJ�a� Lve�龍��T,2�J�F�d���K$��7�4�D�_����y{e3���o�)�F	sա!����5D>	�y����F	MAw�p/�1=��te��|,��yp�� T�����IpS�ΒHiƋ[1��RL��5��ӄ�y���6L�U���e��dt=��cЦXt#pt#`�ʹ���Y�vIJ$�P�v���}g��/!����'ޣQ��\}�>��s��4�~�/�,�?i�I" >5�*0(�5���{���߳ T����v�M�h�޹��uU�s��_Cޫ��ue7��(�����w=�k" J 5:�w �P�' *�)^OO5����ɊQ]���
<J�Jmy]��x?H�BU塞7������(ca�Pd£�c���z����* ʺ'���é^VC�H���ꢛ�Q��:���E=4�I�y��R�i	��+�h�&����-%�jժ�S��M�R��i(?Jձ_h��xBe����I�|����Sʶ���/����KE��R �R���"�J�,����	@����NR*����>�4��A �X�����n�#:V�@g�xA	��]ѷ��s�1�F�K��8��-|��W����������?��?|��?y�o���X�K��pj"�ɻ�0d�+zڢw�F��`m~ �m���{���������ϟ�6�o
,�@I���|�ko��K/^Û���G���F#Vƻb��b�5��sLJ���޵�x��w�_<£G_�G���N	�W��*�C~Β�e���_>���'Qsv?b�b`e�y��^�0�i�����w���q�ݗ���l ���N���k!�x/@g�9ho:�-�3v�A��������MV TI�B@J$dI~�r8@�g[am�F�Kބ�	�8l5�{,�����b�i��}bO��_�j��XG	��D[��Ȟ�t�������ep��FXu\˂�@ �S ���;��@%��@�$�2U ��|�Fh�\%2Tg�<����C��גEH�hﲔ��u����6�ۂ��)�)vqlm���	��~0��})��W�<�	�����ica�	��AH��Ft|<==���E DlP4qA�
@��;ܭ��N��`�bn�up23�K�ի`����~^�(+)E��=�p����|��8v���K���7`�b�Ne5֮6�ņM�"���!�`oy{!?#�G���^��?��Jxn��2�� BRn��ފj�z�c٢e�?kL�-��q�1b�P�:Ǝ�c1i�HL7��]̘1Lf��f������HD�$�/9
V�0q2�L��n�.���ø���Iܶ�г���#�D���T�3�T���h	�/���T��q����z�	�Ǯ �@}w+I��� �iX|�C�Y��s3�Cڿ2�]�;�
���V"s�
|6(m^��~
�ƳMdo�����h�є�<��Of!�T�i����h�f��E��<�P ��~�T| ��4��E!�)�_H;RyM&��s�>�e�&h6�s˱"l?]���H>���C�k؎mg�P��q\|�j^�E�Q�,4�1)4��h�&4%#���!���s������0[QaQ�Q��NO��PJ�MU��6�G ����U[�@!+�H:r�ʯ����"�"�7�\��g�����{���ຶ�F���N� *�Evd�2�S�z���#	�eg�$R��7S�������0z�xL�:�g��<�EX�v%<����	S���t!&͚�ѓ�a��	;m�L�Q\�?jz��f 5���=�`�M�Qc	����N�N�ώ��Ng-h��e�*Yy�4����|�	VX-�l�9X�v�,E�tX��H���24N�R �2�>��x=X�,	��~����<~�����{I�t|�j*����'F������w���W�!�"{ӑE�L�HE��TdV�#� *�i��H('�n�FDI$"��;��=V	CvM��c�/��2��1�P�劵Y�O{,O���4k��$�H��zP�	�.XIH]�'�Rg��q�i�#��*t��"G�)u���S-��|B���z	(��f�ĸ}!Ύf0?���t:��O��>,{�� Xf�˱4�e:z	�(z4�$�v�	�	��e�%�ΰ���Ҙư>!L�)
kU�@Fix
����iw�c�����C0ym7��َ�g3ї��M[<��b��tDY���0��kD��z2��+O��d�7��`�s�L֣ѯK�,����W�Ƶ.�`��XP}	���l�ԛ%�t9��fa0�3�`;����Q��OwB�����P?��N&(�^C��aݺB�ڕ�� ��9�	��������B���hx�N�~�߼��~���j��_	�b�	|�8�?�䖿B3��?��d��^�w }��>Ps����	I�+���^y�:�k����)T�~���Ì���d&L���cB���4(P�6�����LB�3j��ܡ��_{�3���u����AQ5����:�u2VT����@��'	�
h� ���5�RƎ������q۱��N���C!��|���	��Y���YR� �P�.�DD�d�V�=�OK\
hʺ@_��ht$
\���y) *@��MQ�Qe�>
�$�U��_�����:�};�xO+�)�Ԭ��۸�s�+����I��$�����te{��c�E��}�@	�"̶�OPN�R�z�_	�U ���n����?�s��	�r������n�i+�#��#\�ն����S�Y^�N/h>���E ���"x���xC��x�p�'���c�zmq�V�j���`F�9���[�}��>ƽ���ާo>��ܽ�4��02j-dl�h쌃��z8C��K�{�#�g�`\����ꍳ���x���%>�jVaI{$ɏ� ?z�^��-�r%���� }����K���4[�\����`�����㛟?�w�~��|��#�������o����#��G<�C|��x��ױ�q�2tf���TǨ7�(�p�3��Ƿ��;8{�,�jv�4�cL0���=U ��<m��t���XXm��U�\���;Q|~�Lk�hO�����/W�f<	�f)X��	&��1�s��,��%�f9�&�@[�g��,����J$ZGhv�n#z(��vs�iXf�,�M�ª�C� &r+��P�+\I�L�[ ԡ��y+	��s}
t���͠��*��S-�@e�@5�Fե �H|3��J ����H�VF�	�JY��H�T�싥���8�ZIM�}�W���1H�����UpN�C�Y��w��_�~1�8v����6g8�9�B����k�akj[��)�鶉�(0J��d���Ju㲓�5��-�����E?l۶���6~�����p�<Bc0w�b�7Æ����3`gmO�D|D$rSӐO����won'7n#�9����E[��9��1�%����X�܋���H́����n��y�0�<̜6S'M�̩S0}��5�FƜ��>c���Q�1c�,,۸��v���V�X�����Vb����`,��������Em��@{�>�<���^@�r�{�IY���@C�?� ϪxU�*R@��7T$˭�[����r�)S���b�$@#�� O�]�`�x@-Ra�E�,�$|�� ��-,�JF\Ɏ�V����P_ıMdm�é�uh�v<�L�Y'��IM?��T>p����iH8���cI���i7d��0�H���Sj���"3���P�(��Y�����%'�FːWW���2��݋C��P�rv_܃�����������1-�?����D>#jI��0�����F���<�d�V�P�4�\������1n��H 7��}0���U�������aʚ�9�+���Ӻ�� -t2~��7m=mhhK�F�$l�諒	ɸN�)�ں�Pc#h��BS_=���a��E��
GB^6��#�p�
L�9��O�L��֙a��=}Ơ�#0d�(>c�O�~1~�̘;��:��ô��0x� ��}�F�>�a������s H@������� ��'�v��H m��z����>;e8LV����r�����C�Hi�ETM
�C;>^��x�󻓰X񄊇Y�i�"M�o%����:��)�
�IBP��X�5���k(�v���
oV;�p���]H��ĊX��CΞ4l��}���+9���ݓ�l*�����DĔ�=J��$�JF2�.�g�/�s}a��M)�ؘ���N0�;c]�2�k����LBg�V�W�\%�*cG���\�u��<W��wźJ���������M��aWg�����{m3�^�oƤ�D&���Aۛ�&I��O��w<Fl3ݎQPQWۯH���xJ�Nc��]ԡa�}:�%�n�H%����4�Qڕr_B�sYy1�{���п>��c��|D��!�ש)mB�y6�M�У$[��}���P�Ki�!ו)Q(��S�]�8חs�1�CC\���˔,]����4����ϳ��������{�{F�� ���N<�0�q��.����a��v�����DCy<�j%?�ߍ�(x�(��~'�]���^V��ɜ�B~-������L%�N|?��.]���G����(�u�Ƿc��t�f��|"t/�C�Һ�J�T]�gdZm���H@���Gp�y[e�V�x�5x-:����Y�O'��M� �A(�$ �{�퉿�c�x��Wk�;I����y��;���um�m��P����ȿ����t�4xMO�$AM����:�U T�u�|JlC)U� XJX�L7���I�g�-��J&ie*J2I�dYC����۟x;���(?�R�FϽ�:և�M�T�S�5'j)I$�o���٪%ɀ6X/�L]��@�Q]$� �!�ˑ0t嶮,;���z�O���
����~���~o��uB����f�'��R���<�!^�J7E�	�mw�"�Uˬ{~�+:H5wx@GBhwy�}�+���kvR��:@���<V�j��-��:��?J{�;t�Z].TzÀ���������1w�+@�Ki�:�;���;�ѫ�	��l�;��CVb}q rN������뿾�Ǐ>Ł+p+�����D�L+t��r;_�����`��@���1��0j��nd�U������_�C|�{߾���{�>y�|q}�>y� �����[��h�u�j7�CL�?n��3��:��3<hX���'^k���������G�p��x��3���a��R���۰�� u/Aju*��¨����c�0&b-�̇u�'��y?��-�~���2�Cm梟�|��2A_��0��󉘟h��@��{�v�܋��7)�S[��CI�;�H(�$�����曭�1��ɛ�:v#�G�b~�2��1���X��f�fOMt�"L:�u��#�u�ؔz�zE���:-���gC5�$�42��F 54ւ�a{tԙ���&x��s���+} ^���\�"�E�A��.e�p%��m���@8���`��aT]/rަJF�NNԼnG��E6�N�boX\�h����Wl���qM銭&�me)�i�
�F���)����/�#�Rw�APK���63���v��~�=&��8���U�����{\�X1ޑ>�9Y�=��������G�W(��	1�.𴴁�FK�n������e�MV𲲅7��e����N�%�ml��� /WW�ff�DS#�_����}���;N]����"Dť���&�Vb�2���'݃�e�	?{o�q99,�ް6�B�q��h8v	iip��W(a.8�,����)a�N������r�Z,X���/�:��4y*&O���y�8e"F��A��#���~1uf���e�+��aL�,`�r��Y9m,����d�:h���fC�$䒛��)KQBS�r�d�_u$����Es������.�Y�{n���E�l-�=!�%��V��l#$V#���p}"*�P�-ܧ� [ �-������T{Xf9±@�Ӌ�����%�"W�nqQ �E<�%�p-��O����eaH)����GU �N � �
�
�f��@��t@��Ќ��ٔ��Bh�x���+��w�Y���\�
��L�۬@��%�n9^���"��"�Zvr�];���Pq�R�q�XROHȯd�Uht3�J�R+T T�P5t�<�H�E��"��T(T&�8H�9BH:�*�@�D#�P��pW��,h�O���y=1��9|j7�L���<:�A]B;������pid�.��a���C�N�����w������]���X�:)Z�if/]�ac�b�E�st�¥�1H@s�d��0	�ǌ��i30e�lL�>S�?e��r���4� �� :��NY7u�TL�3�F�Q7�������@��!t��A�P�����eЁ�/;��8�7o\�5.k��~	�9��.��5�oN �!�G�S���]�+RçJ�!����,K�t�����것�kŻ-*j����T���@��$$o�GZ9��,�PY���w$#���A���ʇ4qWB
������,R]`. �⤂P5�R��u�5��P���U���u"��f;�*�Ǫ-�XULX-%�ns�#�Cap�!�}!A�J`s���C�=i�"DJ��n�h�@�	��	�ݛ� hKm��<���� �u�� ���5�1l@��"�i��QM$z|F�������u>�`��l� �D�SB��5�A�t,�hl����Hp1&�J)�.�N�۞��*� ��M�O���A�d�ia$9���ytNc`Lh6�an��ߓ �K��!�h4( jH����?�՝�J9z�IE�� 4� ����l}+�^؇m��p��Ӹ��K�◯��ٌp2˧ ���?5����?���޸����Qy�$���bñLlJA�3�Ҡs1��S�#�'�{F��@�f ��u) *�KB�S �k-�پ5��~����h��=ؖׯ��o�-%�َ׼-�<���相?��^���A�%��M��(�D3��O����>�������-%����lg2͐LG��e���S@T����߁�g���C��=��=a��:և�M-Cg����)�b�̵-��:��F<�堄��ZIh�^M4�,��z� i8��ד�ix$��3�GB)�km$���r��{�?:R2�fG�F�ڗ �����~?Em$�m�:ɔ)�HeZ�C��L}��n�J�-a�������C�{�}Wu4�	��H?B*��Ӄ�Z(:U:����Z�N��{�*�`�m��W�੽��z4	���^�-s��'t���83L� �Ӆ0����q���#=�cq�z�B?!0���e8o�P������,�-��7oB7U���R쉉��]���4���8cH��{��0��|����ITQ�/F��=(�߅ҦJl;Q�mǫ��*>�v[��m�Z�A� S�2G���d��;"�|0�eQ0��æ{�m�Rr%H^���8��@��l>/#�`3��k;K�M�<����cj��Ư�p~CV���4�f��/�P��_��*OVcU�%Z��@�E��I�,F����8K�]�����]`����@$�OF��h�����:BP+B�e�-,rm�!�
�,5	]�%!��:���0d�Pt����@5��K�i��T�F�D(� ��<��9���o5f�.MS`I[ ���=\��U���%�
\z�$(��t�\	�����	�}��* �81Q��+����6%�yAmh����W@Sle�ȣ�Y�(��(�˲=�6Zd������o�$.���D�.�O�F#��8P�XP��T���9����E�	�1j�hlr�@P\0�Sb����@�� ���?G_�l���zK8��X���<���̂0j;�Y����.V6p&�:��)c9�ll�b� oDED`��]���[���?�p?�|��W��.Ĳū1}�,L;Kg/���;R�R�������w�%�z!>&G�6�؉�(��DTbl�ܰ`�r�5�g���EK��`w~�k[{'�,��?�ǧf͞�i�M��=r8�������8z0�M��3�c���X�cS/LY:FF�����Eۣ�A,tX���;��T� h����͈k�P��I$�@=�>Px�����.��$�
������������s+}W6�)���;�7�%2- ^T�O�"�Z�9�������i -~�ޥ^��5iE18s�mRi���`UCh��Ld��R��&�NC�	�|hF4$ �Fn$�O#��T 4�T)r��(�O5�*R�i�e@O���d
�J�s���)[v���!h=*.�A�x@�����ͨ��V�1�2w$$��%��r<i���� $pv\�A���F><��y}1i���}j�mk���:)�M}C��)���d��ٛtq�x�Yk�S���ܕ+�qu��iS1|��S�p�
�ZX��l+>��3�!��4�.��_ �=a�슀�HD'�`���Z��&&ҩ;i<�͞�I3�b��1w6f/�K�5���	�1|�(t��=�@���2VT�H�iBO���s�i�繬���`���X�1�f!V�·4����RR�e#�*!�2��i�� �{#�R�ve,h�U�#U\Bo-�I^���;b��НIHݞ��]��ݓ����Ve#��qeВh�m�G�N)˰�J<9�̍���� jJ�TC��,��ҝ�6�k��(˕l�+D���	�6*�ܢ�����XY$ ꊕe�X]�Ocʱ)g���mv��Xe�ɀۻ1	=�͘���X*a3��(�@m��� ��yⅡA)��	|��CG<uQ
��EC�ƣ����=��j�Ѿ��4�G^�C_	��ic�׆��� �
E-!T��D�>a�4�<yl�O�M=��>�y��nc,�-��� ���0�r��b���� &t�&�	*񜏅@�1������/ǒ�1$pv>.��D���M���|��G���sg�]û�~���E�/��{���P�g��|��{4]=��gjQt�AW�b��L�$���p�{V���6�}6h��'U *��2o�ZZ�W��Y-������%��A�� ֡�ׯ=����U�c��V���'b��1\&���}c���A����7T�r)����R	s�*ohKiR�P��p�2�-% ��:���%p�׳��=�O��Ȅ�jG�l�����	@[K��>@�!�)�N<�f��P�OB�D=�
�{�C�+ �}ty��z�3�ԩ�$6>��4��Ш���Qe��gf�/Z4�t��"�p�VX�Cs��(�Xm.k�hTɲ�ӫ�빮��@ɲ]�:n�F�?4���c�7��:m����mq�.m�2и�+�.z�r�Y����=�o�������vh�;���z�Њ^�����b-�n�/�j7c�H:���a���o1�����5�+��U�"W�0j4#����Bt�2A'���pYM�e��n
=�%�Y?����n|ٰ�]�c��z̰_���+1y�RL۴3�Va:5�|Ƭ7A�e��e�T讘����A�z.��Ybj�V�F�|{�o���.'�bM����aK�dw%/�{�ʸJ뙘�0���c��|��F��4Š����}����b",�<���@f}��;�{f?L����|�2���|t�X C����0�2� ݘ��lW�� bW�vF!t{��IGSL͕�^ Զ���V;>�m�6�+c�cE��D�a}�9F,���m�# �q_]B��2���n'�$�� h��}��z	���4����C��JW<�.P�b�k%nK��J  X��T@Ծ�G�NW�;7{@}wG��"RY��BN[o�AT��	������6��;%n��qMi�"hF�%!�^U�KR�U����/����P�* l�j�6��$�@��ibÉ�%�?m+�W4J�D�8��<O�6��sF`������`�*�'}\����'?8�Y<	���[��=�79H�`�����u���3�	��f����r�96�Y��Ͱv�j�=\=��ፈ�(쪬�˯��Ͽ���D?��k��4 "4��/ŔqS�p�"X�Y����V���m��z���n���ὖ�w� �Y���v���f�<uC�������6K+;l0����FL?�ìYs�x�R��h�3CG����Cѽ_Ot��#���
+�v�Ē��h�	���n�x^�4zk�.�[��A�̇[���s�H>��~&�J�m|	�^P� ���$j�O��������ZK����	T T�K����&�c'�S����1�Â �$[2E� �e�#lr]਄��� �^K�iB����q��N�K;�����H��{"�Ǔ	���nd�9�7��N�&�<�LM5�J)�R��C*Y�JOK�2��m��Qr� z�0��ԈʫU�/��2�������p> �E�H\�_��3)��$��"�����Ê��3�bܒ!��dz3�qOI �<;(§~{�I'%!�:*�'!Ԁ *��6�?�M�.@@;?XXYb-t�l>xsN�5�7�*,33�+�'d�Û�����L��0�4߄u�ְr!���s��Xke'__8��! *	YY�L����3��[�e��ŋ0Ǆ�I0�@�^� S�����0r�x�6ƽ�C���%c�$D�dnR]~&���\�ѹz��Y��`��J��.�2�5p�샴�\�5�"���F)�A�qɯdj m�j��O����ͿƩ�EB����J����و�I$lF5���I�1ȪHF.4�";U!�ٻ3�G�̭VhLI�J���#	�ը2�O�Q/��oI;[_�fx��L�4l m��rC��Ҝ`��uR�6��*�����T;�ʰ��L(�<�ʶŊ�X���rl�(��ힰ>��\�4�cD�����2�2K2�B;7��{cz�e�gwQ �Ҕ�.R�V�j�&��`�K��Ԯ�P�[�z=ң�Ц��M�R�@���;_��d�\�F?BK��4>5�+�m�"/�C�Y�0�8WDQIb�x=8�^�fϧ���� AX�q�I�L��y�����[Gc��j����F6�SS �)�`��@6?�?���$%�E�8!t��,8���>�]w�p��E���}<�KR|@�$���J��������ʙ+�B	B��Wh�~��k��BlNa�<8��g3`L�#��/�
@�B�T�/�j���#��Z�����
|6��Pd���,�TK�G�
l��T�ۋ����O���g(�`�xCC(�Wy<��* m��x׎T�f�k���6�@(���&��m�y;�lOГ�1|r���!�Y�ٖ`ٖ�}KI��� T���bi�*�ݴ�j���b{:��lS�O탄���b����A�!���"|�<���4���8�m�-�o@�(�#贍�A�\7��4
���m�3:丢S�;:es[�:����=��v�?��Y�-��NY.h�d�6	֪R��O���1�x.��EX�M�F�	Z�va��瀶A�����s�����	.��vR�m����BEm|o����x���U�I�r�g�_�+��������������(����#��8�E�(+CJ�/b�#p{8�z`N�-����H�Mh��!���>�����ѡp�ςoi�s�`�	��$�!('~i	p�>�I�/-@��\x%󹻙ϵC{�u`'·�!`k6܊S�8���\0+�s"ܱ(���|`����0�lƚ�#,:"~O"w��=;�¬0����OE�U�0�~�[N���8tq����k18n=��T tu�-μq~wW�^��U�� hO�Y��=���n:�����L���!��А�0�nEpY0�%#�)K�)�=A����2Bh�,s�1���VX#�K�Va-���%c�����J�6�Ӊډ�v�=�	��2}^G%����0��Dɀ;�j渚��,��S�Q� ��ӱ4�[�	����7m7��%��mV�4�:� �RBZm�����R�J|T*%�>	��[��+a�	������D�Ų�T�niW�0��������c�C�P	��i	6EbӉ='�8Ķ�Mu�/B��̷Z����a��b8��",����K���nEG��Âp�с��/+7xXr}� ��R����<�aEH\o�M��a.Z�	��Ͱl�
,���V����|<����c���o/?��΋���o����5�ivV�.Y�qc'a��刉IE~~<=aa� �M��%����aǎ*����x���q���x����*�τ�T@�£W7/��7����ȰX̞9������.^��F����=�FL��sh�Ϙw����8
d�6�m0p�@�G���V��I@<9-�T.�����(��}�#�4�{���J�B�+����<+��]�{�.�����v�g�#�P"v%���P��$�r���]�;,�`���@ӊbqV<�ɒq�kZ3����O�"��?�����uI�@�p��2BIF��YN�P)�g=�PP��ڊ�M%Ȩ-�
Qش����u�}e/2	�)�YH?����1�OKBo� *�Ft
|ʯCG�ϕ^����jxn���'oc��? �Gw&�u��S���2����)��e|@c��H�|��0���-�9�342���dm�kVc��U�7o|���j698b�����C�鳸���;w	�{�!63�|�z���a��5��߇�];a��Ի!�� ^���5�� �]�S�����0b��%�J9n�t�6Y�I3gb���ڻ'�v�ag#§.;Y-�42��g�F{ݶxN�z����~�ٛ`��x��!�pk3w$�ߣj*�Ò�N�!��3�ʲ���.�J��!���
�K%�G�?МJ����!�Ʉ�4%7�*i��h6���H$�JQ 4�ˑ�Ϩ�l�|xl��}�'l2ܱI�iO T$�*8u�Y���%HU<�2�(�tM�V��SvX�bI���T,��P��-`�i�E�l�7[��~�p ���&����Q�y4�6�ѵ1��Я>=	�
�>��P��D<���HIFD�3��Ux�\֫�"��>2��.�FÒ�$���2��ש$����n���t&�քCWƄ֪$Ӵhթ��(�3	��
�Fd\����8��OE1�8PPm��x@��S�S�n��"��Ӱ��Cб�F�1�@�'Z4�%k����l���',u&����=��+.�#��߮þ��p��e�U�!U�
�$���= }4�+��O?��+'��Z��V`m}����ә
��OS�3CB��3 T�0�$��`�kӉz��=��))%�O{J�`��(c@B	b���$ ٖ׻��o �����s) ڼo{�O^K�{&��BU!��* %p��I�C�)�M�|�ŤԞ�N͒zMJ�߉�5]J�[kbȩl�ϩ��p���϶lg��fZK`�����=�<Eܷ����K e�n)P�|j�@;<;D���CA�R�����/ ڇ��k�oM$�EA���A��e�����	���X��N�bvu�C��n�'��@�o#���=�	��`l� ��a@���nA��z�(W��@�gt	�F�{����HO�u��O�HƼ�,L�Ĥ0Ǒ	���0,H���`̎������aab8fG��bK���!�a���`Y��Xx�Y{0�.���7N�n�������p�"59���sŮH{�$�� a�p���9c�'�	s���?V���7���^�K_ŝ/����?��|��~�/�^��K|��/x�v*���������g0Y�����_*2e�w������˒��'�?R���！���Ȫލ��(�B���i�������e��ɻ��������rQ;R����1/�{s���>�p?,xAz-���Bg��X�o���Gq��W��;�q�r-�G:���$�q�������D�ΖS���Q��X�{�&����Qz[�����H��}ژA���w5����* ��<G@�R�/�
�⠕0و�+&�� �,�R��P�T��&O�Yfs1�v6�m��%~��'����Q�b�g1� *��^
o�'K7�N§���rݗvJ��T���+�9�ݸ<]	�Rʺ#�S$�΄O�vޓA
�
p�@��:��(§ظ�5�>�G����[D#� i��\��d�����(@Ŧ�q�R��AԾDX�~�d,&��37s�#*����v�p�v��3��B�4�\�;����^�NOkw���;�-	1���:;8���Î d�	;s'XVׯ������"�s���=�.SsX�[#(0%��q��]|��#|��8{�2*�{ ��$\��2N�����X���޳v�-���(�R��P~G�!�p�*���;ܺ��Ұ��a4?wL�>�6�bd�lƫ/�G�$�o� �b�F+L�2��/�~0c���3���{����ݯ+�j�A[�6X�9��z8��T?,�6�*�#S�����Hx��WuܫBඇ�랠g�}�J��%Ӱ4�w�?2����v$�Fhy<�x�C6a�j��
�T{Xe9�G!�Oƀ�#�0
�dhb}*���/(�/�T�d�O�g܉4ĝ� �f � *�NC�cR��C)H�%d6{=qY��#�ʲ �xH�+ �۰�_jҎ�#�����A��'���~���"� �z��q�J�s��' ����QJ���xDe���kN�Ҹ�k�Cc>�e�&�h:ުǩw�!����t��}0dbw��`G��ZѣkW�룳�;%mt鮂OM=h�[�^���;>@E�^�9;bٚUX�|)�J��o�zސ!1�^Y[7,]g��(\��-��S����(�]��(�xy���[�U@wa�����@���������HټY��$��yz���fv�=m�O��1ӧc��9�8s�O��	Ӧc����ѷ��F]d�*aT_u��E:��qt�3���r�X��-�+��8��d%+��R&*��~�$�i�g��J T�;��m��{q�:$�P%"��i��@N�4��yLEv��������IG
�8�f"
�P�|J���$%7nk�*QE
�w$"�J �o��k.;�6�,/X���"���R{A�ӹ�t�S T�t͒	��TѺTG�%|��L&|&۲���$B(�4iS��̱� :7i'K,ζ��B7���bޯ�jc1��6� :�>��	�����6=� ڽ>AQ7�k�J]�Βy�2~�x� ���q�s},�i@J�!�e}J��&��:�Pź2V�Ht���\&�݊1/a��4%<��V�
��=�OM�f m)5�j7�wTr+Yo6%WBe�* �x?yN:T��)pI�LU�}�@��	�ǣ�����t �
�����<]B�K�
]ggBTOB�@��O&��j	2^8�������^�Q'y&W$��TӬ�_�
@�s�
�|�?�+o��Ҧ}ȿ|6�r0�1��<�uJ�z��K�hHBm�g��� ��cяնI � �,%W��LP�\��N5d>K�M��b���Z,d���|]ːfϧ�}�����vl�z"�C)��}�l�z��g�&.�t��� \k�^�&������w#���� ��ھ��K�SAgk�|�~D2>�#�[�����D�}�ϐ@�c�<��[K���Pt��;ن;�T���d���u�6�z�yH�!��m�a��q P�~>�������z`P~ 6T���[x��_�!︻?���w�_��7_�sEB뫑r�	闎#�\#J^�����b�;�b�+�Px�4v�x߼����Þ��P~�2�>|���'?{��^F��o�Ə���ן����Ɨ�������>��~��O?��/>ś���/?���?��op��_q��_q�����E���C|͆��㝯>@IU)
v0O���ս�q���e�Pv ����.�5ф�h;4&:�T��f�<q:�M)n8�������쯈ñ�B���6N�ß������(U}��/�d2�'Ӣ��O��h25���������x�?+�R+��*��?������_~�W?<ăϾć_|�/~|��~�W?���_���~��}�!N�>�3w����ẋ��q�[x��W��_��?A��rLـ�>K1"`�*WGY��N=�����>�n��i�z���A�&��:=<B�z2t��a^�����)����4�2�ґ| �GR�PC�@t$�A�.�DD�ؐEe��,�3�<����b=m��k&�Cw�$�RE�$ɐ� (��Y *!���l�����P��6��#{a��xL�Q�B�e)�Fԧ,e�R�(嶕 �=^QOE��
�߮H�L�!Uqʲ��`��	��%�*{Ӹ��Ocߙ�nP����C;���t,�M�oH�:m��`����['Sf(	lĞR{=�0*�����E�L�aB멚�N�SƁJ)cAŦ'���8��e1�cg��&c��z�SÑ��7o#���~�~�A�O�,���p@�sB\��g�+xY{��֛P��i����p2w���7��	T���}�	��N���x��SAp�s������-ac�_�cَ]8s�
>�\��^��!JvV!.%a���'�aM�tr���&'̝����!#��⎛/���3�����\�������p�X��f-����-]����zSK��8����6Zc�|L�4�ǌ������G����>w�j�A�Nm�}d��_�#+EU%ҦN$����_���J�T��a�d��j�c��Q|>���j��'  O�x@=w�(!��|��4��jQ��%	������u�ὗ�E eM�æt{�ov�����ӡ��En�Gym	��,@]J� ����R?ĕ�!�0�MUh�ěU��WƁ���D�IP���ga0�7qo��*BA�$��^�Y�)�)ЙLI�Pu"�-�P���H9L0%��6�a��JԽv�7�!�>qG���YO6P*V���' �uU�8e����I��NB$�=��q��Fn~u�a����h�ޣ�aԇ�A;�2�C:z��v�B �e��	Z�]V#Ə�:�H����}Upa�P�isfa���Xef
��03����7<�B����=U�߾{��[��G���������'�#� _�v����*++�wt@hrR�".'~ф��\�SV��������݃;�+����~���x9&Κ���f`�B�[��0:��A�޽aL�%L���t��iiD�c���0�d����`��|���M&����Mz�9�Bq%����{Uc��9締������� Z�Ѐ]�����8$�m�H��xhBI,R�')�ϴ])H.'l6���
���H ��� ��>(�lo�j-)�3ݰQBn��� uR<��T��� �&� �lO� ��eM���$+,!�.���)���HM�Ƣk,�u�ڊH�I���h%�",��G��x�f<��%�7�i��T��#������!�� (˞jm��1�Ϙ h���dD���<J<���$�*��F�s�w�/A�An��d<�u£��|���P�"��m��M�JH��x���)�Lj���D<�_H��&)�5($�?C�F9�BJ��T_1���c��J�Q]x�>�<�j#��T:<�oG��l;�W���/?��&�}�dI�b��/�=���SJ.��'���k�^:��s�ur��_�ؘ���2��|�	�z���3 m����2�S$��\+ U T�S�
�F�T�K^[5D�D`��Zn���, �糤�^+u����R'�H�s� � �$0�iP�s�Ç�O{@ū*c=�-�vɹ������yZ�%��z��`�#��`S@����X�;~R��& ����B��5B���R��������A4��>�������ܯ�	?�����E��+�o��'\�}>'(}��[��=%X����u��k-�.�����(��u��P$��RyU˲�[��?S^'�J���O�����%�(FeI:��߂�UI8�#
�hHsGS�.�y�Z�7��p�ڋŁxeGn��J�.�y��f\)
���P�.
�-4'����$�~��y�~�>��]���x�%���x����;x��M���-���Me�+�v�p㕫������m���-���op_y������o㋏��_����P$����O~�?����H`�G|����˷��#������7�������/��Z}��a��:��Y�An��u�X������	���x탻��ш�*�d���:=<B�rt��bA��E� 4� Z��Ȋh$��3�*ɇ	P��JHi��h�V�) �q��g��K Ͱ��>S�6�,��)���i�u��
@U��PBuZh���qG���M�a��̴��%>+X�xh��xo���P�|6K ���	����qߗ��0������@P�M㝰U��XNʜ�4�i�o�%��#�:�r�'�V��A|}*��Rh�J4��o�,�>@<}	�R/�O���$W�<�V��xJw�qY���\�HK;���ٰ�uĈ1�`n�c���l$e��ۛm�x;x#�)��^��E�K0���P¨'����S���u?�@�R^v~p���&7�nt�#AՁ� ��y�<�`mnG[D����/�!gXB]������G��g_�������[wQ��!1X����,�z3kx�`�;,���u`na��`,4Y�AC�c��5ʸPQJZ&�c��Ⅹ��k���4i6�����S�#��U+�a���2p�Ι����x���(-/C�^�Ѧ�:g�ld�EV�f�J2����D�'"�6��u��+ �?��Ǿ`�����!�i �u`�@%	��V����OoC��d@%ב��x?r<a��vG ��`�%�:��}�P�b7�����k�
@��<�G� M`;�(�C����1�~�LŢL�Bx<)S��#�Xb��#�0� h*4���!�`)ӭ��3�p�e��o���	7K �xL	��[i��A�+M��VO(P��|����Bg� �IFBM*�و�����zx���#���K�'i-��04$����H�Ɔ�022���!�k��ul���&������Be���Q�1c�\l��Dlr"6�f������ݰ��QY�}��e&��#����6���YԞ9�#�O)�i�����uXgk��+��/�V�����wT4|�b������[h�c�a����s�gD$�Y�`�)L�m��U�0k�2,X�
�V��Թ�0d�ht��z�F�!aԈ0�M�C'���2�S�a��r�z�a��)�r��z8[�A�* ���Z-�S�L�L�U$���c���\�+#S�����I�T!��H�fi�Kb�dD��V���Xɀ+��	Ҙmq��b	�A�p��Á/�}�첽`��M�P��>C%	��T'*R�til�T�o� �&�V�Е�r��RB�D,N�Ƃ$��&[`n�5Vl���1s$C�먣��ˎ�ˮG�ѓ�~��O�PD� �V���c�LBw�2�JgJ�P��H�S T��c�� t��O`�F�ө
�9��Qs	���$�j	�Gi��k�%�9���XO��u��N5� ,��.�ޮ4ލx�|�.��YmB���P,:�CC�%TXB{	�ʤ�� Y]e��<�t~o���y�%׏��|-�>x����2�~���w�_P5w>�S��m}�÷��|�\��y}f7�a��,t?�	��i�;�����_ �:��H5�����u"u��vT[�+��>*�Y����e����[Y}Jlܿ�C'KE���r���VλZ�سT��x�=	�����)��	|R�j ���K��Q�}Zç�@�-	�=�d��h!�� ��#��`bi= ���_���|�)���C|�����)^�_��֥�-PK����/���o��_x���O|��C|�� <@ÿC���������~�	����"��m?����g��#|�������߲ͯ�'|'�?�~����u��ᯟ��>��?}�G|�Ç����K8P^��pTfE���2�ߕ�+%�8��cI�8�>�V�7^�����h�]�vŕ\7\���E>8�㆓�8�����Pi�γ��#�J�����X����؝��o7�����߽����+���[�!��w?y	�&�~�%��������O��O_Q�����	�?������x���,�?� ?���E5���]��������㯟��G����K�{_���������ŭ[�x��)ܸyw�]�{��C���Xa�����z:��T��7�q/|x�^���,�}7NE�J�$!Ҷ�� �dG��W tS�#\�F�����(�&�4��OQ �y�/���|Bg�xA`�i�g�V�ٹ)���1�a	�tV%!������I�I�N
��]<Ӭfb��b,�^��~�9��#
���-���0�7{C��"5���=�Å��{��2w�k��ʋ�,�"1��Y���r�X�o���4%!�
B�!s�������kHW�)�O�γ!�GIT T�T����P[	��\�~J"��m�W���rCS�*S0�i���������ˑ��OWO��l'V���A �1ȍ੔!t��R��	��҄�$�Ef!҇v��?\,y���ԋ�,�P{���?l-]a��v���.Bll,��`��{g~�^�ei�쉠��Wĕ�����^�_}�3�N��_`8.ZSSx��!0 .<�Y��G���ޣ���9�*�p�������8��{�GV^	CiC&gb��ZDG'b�<L�6�f̅��;^x�E���D��a���QP������AəmH�-O6K8E�j ���#�&��$�h�z��Oy��� �>�? ������>��i|�o>��IJ\�-<v�ۤ/�ܱ1��l`���|ޓ��&�%��\�w�P.��z���V/�R@�ʣ��5���@i��CJ�Le�l$� �OW�/F$ J�?�7�
@i�W�&��*Cv��>B�����u܇ z� yǶ��b5�m�Ϋ{�����xB�����q�iO)�&�9�q����!{_�l����	����Յ�~{(���u`��������� F]:������	W_o��?"����d�*�6Y S�M�Z�����0��BΖ2$dm�K`(��K(!*-��-�چgoz_�L���%0:��Ä�9|�d,65���VDg-[� �;oo���! >	�޾p�1��R�Ko�}6�����kl�����.��l`݂Uky��X�~f,2��q�н?�u6���>�u�.]����N�t�ja�̑X�f~a��R"`/��tN��tT�_��g ~0A�*�y��؉l^�g����DLu<�����[Ry,�w&"�2MIB����BQ4��J��$�Hҡm	�)�FTqb�b�}��x���n߫T���#��a���KH�ls�`!S�SD�@�DOQ�gT~�թXI ]�b��Ul�+��I*�肄MX�b��	星j�Y�1�j�<�@��Db(�A��TG %Duc��hzM��>�� �D����vOh3����ֺR]��!T	�%�*�H�B�WR�>A�|�"�I��x@���$�E� TV1^	��^+��'c@i�+ ��-S���`P=�b0��f���xB�i`k���K-xL��'���ait���������Tx].Eڭ*�^8���^�w��/E�Me����*�����?O9g9�g��G���/��Z=\��cISF���l:�Υ(�T�nE2���vh�)����d�� �s
�)P��Q���$�i�g��?H��5e<�
FU�$uܷ�:�꤄�
���i�{���P+�'R2�2�&��B�gT>�*��� �=�c-Q�d���}D�l�Rv��ռO�5|��7 T�mW-@%Lw :V�)�?����us�0�0�L_e>�����x����ɷ��%�|��~�_��9>~�!>��#|����}w?���?x�}�>��߼�W>}o����mEw?~/�
�p�[���������;���6�~�nr7����o��o���Wq񕳸��y����y�^��6ξyW߽���p߻�Q_W�Ԙ dGy��8	����r�p��/m�x�"�����.��MhW��=�Iw�>N��?�"���'PϤ��D���{:�i��o	X���u���ËW���/oㇿ>�����ß����c|��'������������?����3[�O�p���ܔ�6m҆���l˖dY����)�c�1sfN��I�̌�i�3m�����4�����=�s�7}�n����������>>�ǻx����}.?��|��G������^�K��}s�|u�}����<>��w>{�P{
or��{/�q{Nu�uw���b�dv>ێ��h�Y���e��Y���p�lν�/�y�;���<��8`�[����5X�u�6�ܻgp��a4@%��sp[�Re�����l,L�D�h� �7|B����(�pkH����3fڪ����J���v�]�l2=�!���onJp�wF y/�US��/P�t�$~� z�=��������=*^P�_B��h���B��I-�Q��
��^�'�F!|s4���%�*��Ac=���O�^�oQ�"�� ��^������0�ae�x�v���!f�g�0����؞Ş��%��l��ӝ��p�e�t�x>@(ϓ$D'm��"B��>�o�<�z.��ݐQ����j�e�A����`�`�ü��m�� B/�!!t�!̀ls򒊐�OCt(m� ������r	���7���^*������77�*���A�����!VE#8�p�{L4�X$dd����N��{�|�~��~�-��:������X���.ʀ���-^���[n�6�)s�zy�#�vtU��	���څ�x\��Y�9O<��k��Mx�����K����w�7�;C���)��Hl �wf@/�,���E�,�;�+��,+mQ�Hh$[���m#d6�3|�$�Lˢ������X� �)���(ATm������p���%�6	.�iX
��K%|W�R Է,���,Á,�,üf`eBX�#�T��r3��[Bp�/&!��%��g�'���)0�X�% M$���/h�
d0=��Ɓ�@�S���֓IS. �7P��G� �!�f�,@�ü;�@�:S�
c�J��'�=��b4?ׂ�}�p�v��O]��7���I#0|<&i��[�[��B(�B�c=�gN�wP �;� ���k���
�@?8z�!=?�%ο�
�rJX�d��K�F�.n2��V_}4�޸	v�A���E��g�@�����b���Z�k���6a�u7Q�ގ��H+�B|^!B���`epS�'2^^��_n��������!1&Bjֺ�c���9�b��+�n؀�������F𜊙3�cꔉ�8��L�2��9+��&�0a[����
�Ʋ��/���@e�xe��}��_���rx ��8އ���L�I��$	Qj�	��)
�&6㊌PBjU��	\ �.6�Pʎ����he�h�hTE�
Y����܂�dD޹a� �:g���~Pj#����~��P�O%� h�V@�����ƎZjv�b����������i��f[<�⌅š���dw�2�6�}�7�@O�4�ZeLhfD�@�̞X��5$W���9]YO�B	�"��ޚF�x@��x/�h��[-�qo�gnݙ����3^��E����i�фKM	���+�2���+!��|H���$C��{��`��<�b:W������i��-	�$#�5A�J T��k�%xZ�N�T�_�F}vW<��� �x5�N4��H/���/D4�~�/�B�,�.[�?�ܯxm�sЛkI�dP�z��s(?ҍ��۰io%ړ��20^�����_��΋p)�y� �E�������Q�m;A�em�#�;�E�z+�(Ɇ4�zZ �r�s����	���컚��-��x�W96��' (IF^&%���$鐒xH�� *�#|��� h��e��>�9\��s�e٨R�J���ƣEj4�s�7_��e�~��?��/���+�����h�-g��q��\/��4*�Еi��ӭ�<ބ�(=X�J+޿�vG5rʐ%I{�hw�R�i_ �+IͩHiJEFs:
:rQ�W���"��桶�[:�Qے���B���qw5�*Q�%9q��5a�&Ƿ��(���l����Z-^c��rC�.���pv0���dA$N��8��㹄҂��W� ���8G���a�����߀�D��٣3�m�N�5����Q�ص��N��yO
�3P��X�S���2v#�9�͙�oL��&�U�sjL�#,KԎ�DS�D�?,P!";zBrJu4b
Ba�	@fM4��RIC���er�O���=��	'�:�E,C@�-2���?\��?<��?:�W�=�s�Buo!|�;�ߏ���3z��u��c]���q���0��n���(c@o�[��c��3��q�b~�+�k�����#�_�(BYL]\���L%�k�z�k�/�=`�C�m����LO�g?���^�p����1V�1y�XL�2�����s��cx��qܷ�A�&)�peh!4��Z Է$� A�V�C�����ݡ2>� H�=��<�sP~�OQ 4X �RU����ľ4$�f��[��J�0�� ��92��`����H�>��ݬxG��܋�>�oe) *a���<W���bFBwR�
���-��ǽK�2�U�#)5[�lEFb4��a�a����(�"u���a�~َ��#6��6faZC�?�0��꫆��?m<���/Bm�>цT�;��"�n�񄍃ly܉P�F��Flb&��ʐYX���h�H��BS{.��:>��[�<���+B����jm���6%-����8�s�O+P*�q�ҲP\�� �����Ԝ|����P\V��_}�������QQ���~�OV����,-��~Eo��&���N�a'm�h)u߁ h�����@�� �,�p	�4���QwE M�LGZo�����lɀ�R<����h�7�e|���U����E�-b� �!�"�a�dYe��UD(Д��c@�.�L��$��y ��'	�be�=�4��� �DS[��������y@���. ʂ) *T���F0�*D��J�ަtB���5����K� ��4%�SLo"4���L�w��y���:�M.��(>�h����B�M��$�f"�?�'��nC,�y��̻�>�`��al�FÚ�5~�8L�8�'O����l�F����_p XR��l�J,_�
�a�0&�Ü����l߿�M[��wh���)^J���8>�k���>����"D"	��<���VI@������PD���&��o�<{�%�ͩ��$Bm��&���<~!p	�3��#���2�P���7�j=��^�X��Lu���l�\K ��`n��V��d���N�2�Xc���j}5nz�&�r[����X�^��H蒰�HB"�+�dױ�S�,�"�%4���mlTD\����dݲm�g`c'����2�!�`����,��ǆ�V����eS�f��
�&o�6��ZcV 4�.�8��8;��j�"���<�	�FV��~�U�}�"6�y�@=Ӄ�C�ÓƉk߫�U �vi~ؔ�M)�����T_��ꃵ\�&��L"�R+\�.Xfr� �L�Xg�g���T��s9�Z��y��s����{�'���	���x=Amz_,f��p��d���r���S4��p������^�S�|N���R�DD��	�1 t,0*��I�q��g	ɵ&4X��&0X�p����w�������D��M��A4by\�l
l�܂V�55����n�2��X�$�=ɘ�� +��)�Ř`%�OJ2��y�K�܊y/���Ӆ��P:!9F�tt������k!��&(a��y,'�N���-�s�M�:P��c�(d[t�����WK؟���_�a�G����[��/�� U �����aۑH9���xzO>n;����3`�?V������t� ���^�qJ"�a�FEC/��t*��g(�R<���M���LY
0�#\0��r�%���F��'��I�/�ʡ�D��S@Q�^��\I��x?E��|�R�� �\k�����L
$�Ww�n����
8*�1.e�SB��]���֝��+��1�+��zt��+�S>�����=�w�J2�����I�l�oa}���r9���Ԩ6�r��W�i����5<�� h�J�>�0�!㛴���{2�Q��!|���K|�7�{u��  W�5)^X����x*��';��dG�Iu�&����o�}ԝ���Ǹ�u���ո;j=�6l�~J�wG,�]��q��\<�=k�V�#�	�,��k��Y��Xl�jBSK
��R�e�[�Qݚ����PTb@vj(��#�W����I�K�<H��Tie��X�Δ��L�'	
'+�8Ueĩ
�(�����<��3��x���2�*v�z�����[u��5��^�m��Ж`�Bi+��V��U���iz[�����ⱍ�qۊ;p��{1sý���aL�x?&��W߅����[0j�M��vLY{?f��=��1��x��I�vzs=����E���0� ��Eo�w�+���4&v��'Ņ g[ޓߋ-߇C�&�����P%>��Y���q�}i���O�ρ�z#T�j���`�jVx,A��m��������CpOU��:קp}�"e�+�G`e3O���eC��!Ӈ��E �y@��f��Ӧ�4C���p�T�¡HƁz�.��э��펍)�pN����K1d�P�3� 9Fq$���1�hB�d�1f�"%��#�����Q�q@X����ci���I�qݽ�a��'��S�m;w����Ѓ���̑RFۮ� ��XJ0 \�E(
)W_���V�%��i��(���J��Т ������i��
�����¹8�@��g�I�YI(D��K#�%�VM �Hf[J�0�h�Z�9��ψ-狀Q�ߊmE�l�%����@c�hSue"�#����p\��V��ZhB������\�#����*H�p*�?*�0��|C��p�`E^�sW)cF5��u_>'���\	���t�gy�#hn�V��hc&�|����^��$�j�cʄ>6AЀ�H�S���g���e����a��ց��M�>@���=��G�@�GX��U��߱�O�!pf��v����ҚZSR���~�p���лs'^|����;x��7��������W�8s���	�fM�=C��3NK�ƺ��_���td)!����LQBo51�h'��@[�i�)�q����]�)�9v+�O�JF\�/ǃ��E�`*�VEP!(�ߒ���|�Zf@@^����'7\���.�|�p@�@Yn�&zK�,�O�0�rL�"|V��Sa�*��6����֞���=CO�4y;�A�;2M$tJ欄�4���]�9VR3KV�(ť���X���%�'�sB��x�@1�I�ϔ�\��"����7���n��G*sJw"�v� ��i ,�'#�/	��	`Bd�������"���d�O�F�]I�o�A\++igA)�{���J����Y�w̙�	3�����l�&����&b��	��崩�1l�5�u�,�z�����dƢE���s u�yY�)·1)�x6�i	�N�G�!jC�2ߧ1��R��LfDĚ��BI�II�*�U0��|���PS,��b�q�q,�1	I��J���,�x�v�+����ҳ���;�<���N�apV�1�"&~Q	p��{��*O,�`k�t%���E�c�M�1v�5&^;	�gN���j��1n�X<�ԃp�w���l�l�ܞ�\�fKB�m�T�Xp�+�b@�Q/s�05[%�&B���N'i÷���"	���"���eB�<$�)�m�u��xu]�i ����\����nN@Z]�M�.�+�}��P0U��\cR��4$b	��?�*NYY	�ب�s���G�#f�Ng�L�w&A�r��SF 아D~�O�zj lS�a�쏍Ʉ�?l���d_�I���Bh�V%yb%+��7,5�`IA�Z��4���[�-J����*��y����}wo
�؝���%�b	���D���k.	t�lӺ~[ʾ�1����L�'ӵ�$0�g��\��.N�K�8�¥xbd���-X7kp��$�9����d�N��[�	|�`k��T<_$��x/S�{��ޏ��L	#cOe:���q�n_f�J�u'���G��f��Pf������h6n M�3�iY�|r�^��	�I��);0u�$l2��b�T�aG7�|`�u�O>�ϤM�_�W���- �G�O���τl�����NCށ6���b�v>�=��u0�$��`��	�&�[$�z����pgP��.��?�g�2	�]Iz�e�u9�{W�J�;��`��J<���(�3(�=��W����=�!]j�
�vZ��]�x(��+�
0�{2)Yթ�Lsb��0��}2]�UXldl^ŋ����/�d��������f�Hj���4nƈZy�f�6~���'��x?	��[՗�~�f�Q[B1�>㷪0:Ǖ ���N�+��O����C4�ª/��	��m1!n-FŬ�И�:~%�%���������(.G$����5�n���;L���Du�&�rݼ�#����1G� �7"&_�rBf[ov����;�L�ۓ�=f��f¡�t��+:3�����Aq���#��X��ya8����8Y�����lq(N�ip�ʀ3[�p�!��ൎ"��Q����8Zm��|����)�uQk���Y{Ik�%z��mё��˶X4��`+��F�y�Ȋ�C��K���6�٘��(ƸߏQ^c��C�� F;=�)>�0��I��}�0%d%�Y�"7b������UxR���G?�k�n����}���-
���p��rM�l�a����߻)�c�Qԑ��:��^>��_:����@}g)�����G���;F`��X������/���'�w�~�*ܴ�!��47,��ʽ��t?氯s*���lo�e����A��o&(��bc��'O�E#���Ԇ�|?8����R��BOl�s��,G�|	t��@�°�C1f�hXM��x6)Y�4+#��+�y?Gr߈q�1��/�R��}�HL�2֓�Лf߄yv��<���.�p�����h�*��0h����$a:�(Ań˒����N�)U!�
�sɺ�,Q<�@��+��y��)��o�/%��C�E�ET��=f��i�� hҶ���+�%� ���)�?H[�fJX�`4�`��zZ�n	;[\7:�^��D̬,��L��@��Jۉ�=��i�;&�������M��@��d����X3���Ѵᵄ��0h��	�AN?Dz!����':o�˞�U��Q�.���J����w�胵�`�J����WG�0�;<��Ժ5ې�]�]��}�*5"���tzj4"�c�iw�;���Vf�x�����W���W��+S*z��!6)}{v!��U[���qd���)�Ԩ�HG�^C�յUx����o��[�q��H�O���Y�'S���-�W�>���6+iO��8����$h�;ڻ��U��ÚĔ��7�����Qn�DhS�rL���x�z��u�P@��Z��j¨$#�j"R������7�WJ�l�r"h�É��x7l"���=�-	Q�������SN۸B��J�eBgH5�5��J�z���\���X�ǰm��@�9@���.���,�DEQ�,���)�zD�����*a����@� h��b��Gj;՚�ܮR�hD׹^ԟآ hR�)4X�� �xH/��VD#��ܕ���T$�� �?[�m@����xd��w�5��2�\�qcGc�x=	����4i�ej�I�a���}(�*���+��m��D +'��H�a <�����`hb����
�Ɉ�HRr���������gd!6-^a����DR�UQ)�������L�R��DDc�;g7�����A1L�� 5֮�������cC�6 Dk�w��������jWoxG�੉��8�ã����Ǘ��3�6`�F�Yo� �C�h�̼e��0gY t��фЫ0�	Xm�
ؤ�5ZrgL��B6l�J��+����CBf#��s)�ϋ�)��j�
�J�R7ʀw©r� �N'����'q4$.�A	�J��j��	�	�4,	ձ0.�L� l�K�)�U��q�q
|��y,���"RC)��Xm���:���b�z��1��4��_P��+ܱ��e����&W,�w��Ge}�����X����z,�M���T�Z�Ƭ�p���s�@n�iX�L����τY�q��������\�B	�<gf¿�>�(�c*��̰&$���2_� �U������N��{3q��@�0�yc:d
��X t|��x�dދ �X��S�MEze��t�� ��3�������;�% ߴ+7>��eƵ{0}�w�t-xB�e�PB�L3�=�ЫS t��4���"nO-N��￻�;H8�� @�S������7_E��V�	�w�]阱7�Ot$��$�Q�ԟç���i��������{����������|�w˽Z�x��xOW��5�z����(��0߫�5G�!���)R(I�5R���(����Kj+^P�s�ؼ����	���\o���*^W�ܯ��U��!��"^�j�5�0֫��#�#��Ϸ�:-��5F�E<#0��9���Ik	���0k
����l�� h�;�����7�>���?}��y�G�ٞy�n�#n*����U����\����[�A�c�֥W�	e����tL+��|01�3��pc��OوՄM�E�W�vWa׾j��Y��}�8Й�C�-N���m��웞����.�/fO��΃Y�]4�����D�v�z�p�N��T~ �%�!����9�-/lK�Mix�9/Q�k	��ahe{]���+Q����ӮB�~�F�G�a�c6�%ֆ�#|:����H�l4�Cm��V"����ZW�,S-�#*����0E� "a\�bLV/��RL�,�8�RX��c�v�#h�����볣�(%�Ƶy!p���ba_�9XS����������6��	�K���D��2�w����x���q��&��������nǭ��]��t���V �eB3icy,�m���←�����=�'ͮp�}���le~Aދ�5є� K �W"a4��"�^׊@���Ù �T��Bw�Q�%~��a�j-��nĿ��o$�"Y�}#0FƀN�)V��6
7?t3��y����qwm|K��!��@P���B����@I�_<�O��.��l�	�
t*"�*�l[��A� �;�>�sʷ�W� �FQxM(t$�>NaO{�H[��nI>$^M��M�1�P�W$ :8��2$��^Z�,��F����M���	���6��I�~�ym^7�-Q�,,>\���"�V;��0�v9<#h�������6�u�*ә�u���#���I�T������
� b����l�14��p��7'_x��Ã��[ ��vN��|"i�������X�v�ƞ����WN�L@0m]o�P��a� \��VO��ę��c�>~��U�q��I|E�๗����W-���2�[�����O?FI��g�rr�W^���RĚ̴�����><vϾ�<v�K.�ǽ�oǐd��!�������ܕ���y0��"|���T�~����
d
xFЦV�q)*����ڨ\�l�uB)�T�U2�^<�2s% MjOC�vr���b�mT��v�&ڥvInpg]�-�1���@#�W�P�m�I���+�5P{@/��%m�;GQ�lFDe[��$��+%��jB2�N S �^�?��}Zw�; ��(F��Z�>ہ-'���{�IB2��@Y��(}���<��s���ID���HEbW&2�Q{zv�3���؅�ǌ{�+��c&^��G(�`N�4��e:���&c�I�����
B��
8z�b��yHOOŧ�|��YX?��؉�(�,�!Έ�0��`�tjDD�0���`BAy)*��PXY���$d� ��U�ZQ\߈�-[Yȷ�����%0ed����̂"^3nPiu�4�@o�GJJ��+���ud��;+`��G�ь },�����@c
|����Wu<tqX��g�k����!Xb���,��d��[�������	�&b���5i$�Z_�����vp�q�aJ[���L%����ղ	HFʸM�����) :X����@ػ�,o|׉,�2'm�4��W�H�@ 5J��-�6"�<1EQ�/3* å$R<��@�o�P�e�O��5�F+�Be|hdaTyd�)cA���	���"|ڤ�{ ��'ͥ���agO�]ltP@T��_���?�퟽��Nb}U�����H�ߚ����qs�����x�#���D�r*�e{:AtF�3	~3B	�3�0�s]��(:�׌���^�EK�HL ��$<��o����\&Jcצ�8��4��v�1�ǀq�2�(A���ۡS&��s$�W T<�J"$�3���۳���>� 9�טJ���#VIF4��hJ�f�̸2�8Xޯ\cFO4��aª}�'���m����_$��o������_}����;��{J���x�1^��j��?x@T S	��|�~�A	�]I��!���?��oPW:��$`(�C��8��W����r B ]�� �PWc9�e_d�PD*���Ep)!��N�O?���1�:��9����'�/���>~��އ��#@��NW^k�|o�F���Ȗ�jU<�0f[(�lŨ�!��͡���M���Q��j��\7ܞ����C|�������.*�w`���%:>}qAw��B�+c���0��CK�0��W�J�pM��WycR]n��)�iy��.ە�ဧr]�Y�4�3[��p)v�bOO�3��Sp��)�g��q�3	'�Ұ�U)>p��0���Ķ��OĮ��V���lϏ�O��d~����D��-��Ж�g�&�T�	�j�p�$��>�����P�U�KQ�^�&��4[�6��AQ�a���>r-�Do�6PkQ�uT�q-�"W�@�&�:hVb^�L�{B�4`�v	�h�`T�B�R/�H�bW-�h�
L�X�����{��p��6�̓���Ͱ���R��*�����B�$�Kr���Z�၅�nx&�O'9`!�YK�j�W���>��	��9���\l�؈e�X�O�/���}�:��_�P �� ��7b^�Z����.�uA�a��F�>������|lJ��g~�|�ћ��VF°ŀ���Jd���������Q��@�
����-��S�7<�/�.kt�~�@%Dw�"��1Pe
�I�\�)#q�����O�a�����v|��FT�	�a(��Mc��6� ��aJd�,}���R���*�)��`�������/&x��'xz�{+X� I�v0�����8$�_6u
|�{��^<�"�|*p�d��xBE�f��ܥ�s,P���h5�4��)�)�Hn�(�H���$�e��L6�i��&+Clq���X�ew�bӓ����/���*��(���D!6� ���X�����!H��bBi�QI�dh���f�wg_xy��# n����A ���=��g�GM}>��;�y�U$g�����h�1�`���3"+�I���
Â%+�УO`��z�&�uѴ��QM�T����Go/��C��]h��Dzi1Ҋ��َ��N=}
�}�pw��]���^8�������O�ؾ]ّ�Ôy?�;�D~k1
wT�cȅI�;�֍���f@8m[��A �@�xEEjB��F�x��'�T�e)�9���W�T�Q�@�@K��Q��Q�-#v	��dr�}�+�[���[oʫ4� �"���	�F@S�ARM<r��н�N 4iPɀ��;�{���7i{(Q�O�z"ϓ4�⥊hd���џ�t6��2�����+ h�$!�*@FW����^��5�N���+�_���=��P�d�LXl�|&))�M4�ӷg#w!�^�BÉZ�x��������P��Ic`=�$���I�4}2�_?7�~3��8�|����*�>,dI��/i��O~��4f�x�u�5�!5#�X"M8b�q(d�����ֶV�:x�N�B}K+�;q�ͷq�܋H/,AJF6+K�z#��P����~4�u 3��ɩ���Q!)%��Ş}'X��������b���w�PMB���3�1,��i���.D�5��u����Xxj1��w�Grv"�xb�|\�M�q�LL�qat"�����4�W=	w�;G�f��ܚ��~�{����X�����O	˕|z?- *sNY T�5����e��2!�P��+�x@��7�_��*���"�J
��U|Z�S<��W
ǵ��eL���DA[�Cx���*x�R
�:��8>eܧ�������eq.XJ�\lt�"���]����4m`+���Wx���,c��xuo��Go9f��n6�V����0��'�9�� G�����O]�3��L��?�$3��uj;9��e�ú�HcW�	zF��	����↞8�6��[�3�G~�$�x� �5Ael��!% H'Ȕ)����R�r� �D�d����'!��<>k{,�s{2?;� 4��i�� �x@�K"B�L3� :�P>��u-?���k��@}� ���y2ջ��<�����J�����E���H<�n{�1g ��J�$��Ͻ�(�ᘝ2�S�^��A|� *a���m��~� ��$��/�ֿ�!j\թ�xM˾߾òm��x�Y�o��^�!��PE�/ :R�� j-|�$�d��]&Z��h����2����X�65��լ3����$3���h~�H��\ݮ�}X~�x^%X�GPJ�!�)�|
|��4C0��9j+!��9�!��=R೙���}���%���]Y~h~�8>������	�Ouc~�;�7�`Z�nf���^� ���	 x�cx��)����W)��5U>��m�#{205�c��?Y  ��IDAT���G�(�Q&S/�m�}� �i�������?g:�q�3/w�८d�a?t�!�i\W�z ��Q�/���M�U��ϞT�:% 3�p4+G3���U���Di�3g�p� z�)ǫ8P��w�iס��Y�5�U�Ӭ%dnBk�:h���9>	����O�:�Z��סް��ը�-Cm�r�D�Ba�r$i�AGԮ��v9n񛃩�s06�)��X�a�ϡ�(�G�HC�al�
L�n�݉^x8- ��{�&�:���y}�K�ð�8KLˊB�L���xc~�'���\<A�Ou��=�l�����û��x��(�(ĺH,�m�b�F<B��q�[vo��±��xT9z���4n�\�x�T�����m������\ɕ ޕ@hk�C(!ȉ��D5m���ܪ���ep*���/� ����ė�o$�F�c���2��~+��J�"#:��>�/(�@%�œ���I�Ŋ�"T��v�����L�R
_����h�/��fHy�2�S���-�QR�e�e,�oA��-��[��}~J�@hpyB+y��\MCb�c`f�l꥽��9�G����j��VBl)M�Qߩ�%���a ]@���:n˸���z�9����+a��P#�3��6��-Pj[��]"&�{K���y����N�ۧ�Ț�����q�9q�}�
*��/�Q:=�L��JJGbt<b�1*=�C�0�F�sO;5^O����Z���pxx����>~�Qpt���B���ډ�����{	�%U�4��?��w*��e0C�g���hc�C��`��f?�[n����ǟZ���,�h������_�g���YȮ(�֞.�:v�~�%ν�"��9�CG����
��b/ȸ�W�z��:L�5S	�}�釐R������(Gro.�3CV1���LP�ڶ����x?c�|G��xA/��PJBsh��	eY(!�� 4�3Ż�Sk���T�#���e	��@e�#��z@�	��Ph��BuE +W#��ό�lFY<:�7cHJ�@3we!��;k_.2��+��� *�����=M	�5v�8�l�AޮR%ɐ�fҠ����4{G)R;ymhf'����{��}����Ԗ��.3�w���T����X��x�[���>>�}E�|�z>�ys0��I5��I��7
��L��I�0n*t�dL�vf�zn��N�[��]���灊�Z�8�YY8t`?>��S<w�Y\�p�|#�g�����/����'QTT���`4l݂_~-���طee�M" !%� �1�����;<ܽ�����慲�jlߵm�}(��Bbz&�"��D�L��ɯ@Bj.�Y)m\���E@��[P8�B������?c
�S���7]<삵����n�Xe�5�X���*2���w?t?n��6>�k �v�d5ny�Fب6�-��I^���FrO&⤱�l�
BU�y<=��-��ؔƏ�(��,^R�Vӈ�.�zd,�V�� *c@U�j%	� hS%?[��R#�j̈�$DT�����{B4���YB�$�ʺ��)c@uEzDHեz�e����S�o �1��P�Vƻb9As)�s��A�%\�\L}2|-��� ���Р{秿�+6h2i���	�͸?3����e�zvB3	�Sۢ�:Bg4�	i�V ���	�3B;%W��I]י�Y�_�X'v�(��V�O��.���4�
����L�]{�q���T�#�7���+����� �8^k"AQ T��ʾI\N��T���L�>�� ��� �5�ŊF����d��I���1��Y��=�u{s�;RǶ���x?8�~�Xп�l�^I���Iv>���_�C��Hٿ�����,ܸ+S�%c� �ʘ\�X��n3�v�+*�P4� �3(���o *�tAI��_�|f:/����iH{8!4�w *Kپ��"��5-�������$e����@�  @�j�z$ \��z � )b]���[���xAy+�K��J��R��j�P�gGKH�E�\����[	��ϑ-�Ֆ mİ� o����F�$|o"�H`�%��02��d��� �5~d;����=݃yqn��S�#ʽ1�6#�<1��c�}1��CK	�E��g.�0��c��0����q��+��#Q�Bc�7{{Rp�=�:�p�7��I�����4��ј>K{e��P������f[!`�h��^�]l��	�����c4��d�)^�cyAxaK<η$�x�'	G�ؿ.�`{�asJ@��Z��fWt$z�;��i��K�CW��PKXk4أ)�[�m�kQo\������.Fu�Tj�4r)�5K�j*@��Kp{Г��F�>���1L�W�.�5!02d1FB�bb�J���d^~8VV0��kQV0VD`ea8֔h����T�a~A ���œ��x2��g��t¨#��ZG�-��&>��E<waμv�pL�d�e��Mx��`e�z����W* z��C
�ްj��+c@'y��X�9����R�)�k�� ]��&���#���X�2�QBp%	����W�U�g��
<`G ud9��s��
ktvu۸@	�c	�E]���0~�Xϰ�]Oރ�����q�<�e�1��%Z�����'4@�B�MC�Д�BA��f�.S]R	�ɱ�����3@�T�
(��^
��V#�*TР�@��D�����m���b3��ח-�m2��2��d�O?�B�L�"�I0#��L/���[�z*c?i���OY�dD
���.�{=�v7��;6��TB�"�!t��y��g�`�q��(�Z���Ź���B�9��)0D���@C��Z��NMH$bh�&Ƨ���)��8�*=h�J�w�x��B��Q���;�k�1T�7#-�}<��|d��#4����H�{#TE�SG_<�4����xr�<��2�^k� ��~� :ތ��r�,������ۯ���l�GvY��
��ן�?|�_~������d������1d�U�~׵P%�P��{P��:��ā,zd�O>��%�m_E�%�A�m�T�S�����Cr����� ���o� 4�-�{*`nLFx��eP�$���	&��@h�:�9�>%�P?����S�� ���ZƀV�"�Ѐ��JI�T��Y���M��ޟ�@� |J�������d%W�au��h��,Q2�
d&wZ��L�ɳ��^P��%�D-c@%UzJ�%	Q���}[�����r�i])J��)0og!@��	�}��O)���Cg�V�HR�y7����xk���B㻓�ܛ��]9�z�廋���mO^��G`��!�0e,&N�q��a<�S��7c&�#h]���<3�<��@|N*2�
gDHH�24,,*TWW⣏>��~��{���9>r۷�!7/q�xDDF".!���/����;��܊8#a�H(O΀*$�NncHL�P<��(��AݶV��:���R�Rr��K���'�2z���/T�PG�`�{�54
N!:��3��,$|�a�{ �cRᩉ�z��_逕�<��@�+�1&%`��u�c�ݸ���p�]�c�a5m$�L��vs�nt���A��;��Yl�R���@x�$��x>-Yq-�p-�A�$I@$�n��|l\c�O�H@T<�z+b8����h�u����X� ��i�1���زe���=:/y@e�hi4t���*�D���adc* ]��KhԎ�mK���$�b��6$�b=�sM�7�<-��&w>��%4RFe}y���܄�BV#�6g�y��{�_=��?{�~��F����ɻ��1��7C S`��9U��-:L�d�LB�t��$<vJ�SY�D�:�0�ט�-���	p	�&���0�7��h	�U�54pG6��(������������9��߄�MjLl�( 9�WEB��G�O��+���O�!x\C��$�RNj"�O$�N�9�x��;N1��XJ�o�����`�d����<���ň>R�2Z�}��R\	6�������{���c�wU��lܺ3�L�D	Õ�@w$�zG"��@���HBq��.��?:����� ���5 �H-c>%��G���;�^ӥU����s���py9�^~�U
��⅌�P��0���*b�N��T���Y�%��cFnW<�ʱ�ǯb=��-s��oS�y�uG	t�=���&H@�$��a|��K-��]V-�O����K�$��$|����rȶ`i�2 C�B�_���wU�?�4�PÚ�0�� Y��`L.���l+O��_�ç��~���<�[0��#+|0��0<����1<��ݕ}���|W�u��,g��rí)�x$�	3��+�@ICZ����-�v&�B{".�X~�}���k��q@G*U�Q�޲�o3�(�+�O��G�#+t5�WŠ?'��������6�(A�8�DN0O�D��3η���fU�p�\�]�A�j�E)m�&�Z�N�J���_�lľ�(�b�sї�ά 4�xb[���fg�F�E%�J��+	����P�Y���EH��h�'�46�����qm����rx�B� t���?�qa+`��=�c��|L
[��c�H�7����8�	�K	9�%� K�C���4���x�/�ǲ�-(�Ó|�G�D\}����/��oǅ�N��`�2�6�U�F��%p x��n��E��Wo��+G����ĝ>�q��"(!�:t�ݘ��˴J�߭�-�Ʉ���؏g�f wo�bש�hxw���*.e� -�V�9>m��
�n08b�m�>Ff4 \N����j<m:��r �$ "d����cFc��1k=V� �ge���Ӭ0f�����x�u���|�k!��-�J�&e
I@$P?>cQ@!��D� ¥?ԟ�Y�%{hq0|��~/�Q��A(�+T Է�F~�7<�=����mo^�[�M 7�İ� �I8;ҡ�0#\��O9���GAE���^Z@U��D�(	�m�}1�V	t�:Coei�ʘP�pA�6��Gf�Ȃ�7����=P
��`�uZ�V��r��tCE[=����>qP�P!4�`�3 RM��� �v�^mP�� S�"T��TB�U:�q;�����uY�d`˶�7u`kk/���������O�&NY�����A!QHL�G�9��Xx���z��/Y�y�Q����W�Ņ�����d�ػ�ۏ�w�ހ.9��b���n��'_��c��~�G�={/��)V>�
.Z/������NaA={W)Rv�)/�k�mhڢ�����{�r��M�����6�� �q�����w'(�$	Q�V�P�7��Gx����/Bl�My�2ԿP�� ��;c}�-�S���b�����|V�lW� Yo���> %�U��H u�Z�Œ^�֞*Iߑ��~
��%�J�� tBe)@�d�m�Cz_�2K���
t�xBe�@1
�T* *!���(��HЪ=u�y'��iB:!%��mRo��(Ӱ8/�]@Yr!T T&�Mb��|j3���1l��nz7>4c�]����x62S�M��g㩅�������ٸ��q��w��9��K�N�
Dp��Q��tp�p�F��,�.������
�q�����[��Oc1����>���>u-��,����ڷ���#.���?���
���yk+�Z:�uk*�k�����>��T���#��u�hE�H&P�RsmJ#4�(�M.��
aa�*ڌPC"B�IЦd#4!v��aQ�u��;ou<ֹ��'s<B���j�a�H��s��p���Dg`�ָ�zn}�؆m�!�'���]JZicW2�Wd�)�C�
��xR� ��^�z����Dt�f~�is��_fPƀ��*�?��?J�Ԩd����<a4�K�����2y�J�C
�3�������6�6ɿi���G ]I ]erê��K��ˌNXㄥ,���<���^؅�s�q��7��g��� |�b�4;�G���A��NBk/���� *@:CBp/���L%�Nk'|@�@g�#�)����e"|�@�
�v ^P	)�Ih�kƨ�LhQ�=�x�X>�%�^�s'7��P=�C�E���BȔ��4��:4�Q,�$P�t2aG	�%��h��	��.zy��AJ���@'u�|���=
����h��"c{-��R;��W����~���P�����x�;7�%`��LR�o����A���ƀB�`�l� �&�&�;@��{% ��o�'�9x��^M]��	$��*^M��%!�J!���ii�����z�,!�k��cY�&��O�d����]2-K&����JعxJ���>�������z�h�f;��I"dJ�N�i�%2a���q��mZ��$��V�����E��uv�,圑[C1� :>�w&���X7���[|��7���/�saŸ���M�Uዑ��bw�($�<�d{h	U�����I)���(S��f�@W�B��4�w8O��}��@�|�%gi�f�p�^�]�����BS�N��c'�q��O����g���t�.����؟�c�a8U��i~ؓ�A ������W��2p�J� �>�\K�����o1Z؞�6��x�@^�U��샶����`��0��;+th"�РkLtCM�T�נ2j�5�J�g9�(��΅�otAs���=�{B`Z�b�W-Ǥ���9Cl�0����[�1�1�o>�{?����a�L����S=�`�f���A�Ku�b���b�&�>�C ��Ƽ|�g�7��t�I�xL����?�7�<�W��|q]'����%ћ��䀧�k����s���#|��p����7�.۹��F�E��3��k�ޅɎs`[A�T��z�B�Y�؆xe�ح�0����~I<�nPIB�\bIB�\�s	@�
�V����C�5T�L�	�JJ`t@e}B@Ǎ�¸��o�I<d�q	��Fc�L{�$ܲ��o�t�������u�!%8��xA@��,:��@}	�������C %�(^P/�x�� ZJ{*�v����n/�˿�Ǭ���gH��dN;+��!�߃�u�D���yg��Q��S$� ���x3�O�h��R�~>eL�2.���k�G$m�H~>��pڛF M!�`%��i���g���X��1a(l����}8t�$��K����C�
�"�vjt$m-�C�^���p󃻛$"�g �h㪣bi0A�{1�kNGRz>��R����<��L�bc�GgI^�G?����F -�ڿ�Z������?l7�F[f�u����
?�Pe�O�N�(�=�8{��Z�I!��:`���1�F+8x�G��f�9> }r$�f���k�b��&�m��s߾�7�!�;���H�%�+�AC�T����Z�s@KP�G �q�2%� ��6���Z�IH�ZP��P�V��К� �x@#��R�g�S�3+�l�m�NpH���z�L������2���\@%+��5��,��=���3�~K ��̽9W�����1�	J�da"�32T48�S�S T�)�ϝ�
�f�sa��Y]%
�V@w��M�nCrG���� 4�G�p%���P܋:�M	�ŗ�{ϧ���7��s��ZZ��;�:�^z;��a�1S������N�Ó��#�F�磦�%5,�)J6�]<C���O��"<6
aQjD���g2�QPZ�(C||����Ct�6n��_~����=M=��|����?������G��k����ӨohBf:+p~1jkp���x��w1�{J+k`NMGbF&b	�a���]��Bni�[�Q\݀��ehvq���%ЛR��K�}'"���$#��0U�y�Q7u#,&Z?������O0Vl��WP(22��9O?���	7�u-��2�&���Gc��x�z�-����kO��BLw*�3Q������
�����Jh��3^Y�6D#�N1�q�bJ%��"�VJ+㑰9�2_
���g�2T�n@5�j��T
��s5J\�4�8J	� uJ��F2	��	�.ş
��E٤`���^@W8��Uq�XN ]m�EQvX���X��ά*Ƿ��|�O~��9mK�({x��6�0�%R	w�!�IMk� 蠦He��6�� �. �:5���"Y�\�T��i|�S	tS�c1���N�������@��):Bh�ڗ�[L��/SZ��5��єqk����q.����'E@ ��3�d�!�1Ǹ	d*��u+��5�+t'IXr�3��x���v��]���^�����(��$4�~�*t��� �t��6�ɳv'c�~kбPYZ�W����P4�@-Ʌ��,!����������?�@�l#p�����c�] :8��nK�CY Ixm7�S��c��-<?��b0��1i^����@����u^ FP�!U���D�b
���-�Jt�D�sk��V{�?�(�HǶ�m�ń&֕jB�\�ȟ��Q44Ƥ��*��Y�����(�[�a\�
�۴�-⒆��cl�
hߛ��gw�;�_����k��:��q���[��[�a%�BW��P�B)p�qM��f;cj�nMr�B�#�X�r�W���!-&n7+�s�6��mrb��iT��9bK�4�w쬏³{Q��9��������a���h�=�>ؑ�}�8Y��%Z�M�F�����js�!��ѓ����.
G_�j5�L��������]��Gp��OC�7Z20P���=�ܑ�D��ˡ�y�>� ����/G�KY�
�k��\�e�Q2ف�#����ρ?�rS�"�[�[B��ڰ՘���u�Ickυf�8�;����� ��<��W��x�����G��#�ݍ)n���Z�#�-�
�¼ ����SY>x,�';���e�崶|�������8{n/.�u���uq�X���ڵXm��}����/��^���!8C��6��M��,��|�c
u��;y?a��`"~�d�4��(Yp�|�q�$z*����55�J���$D���p(�$��Å�O�ϸ��c�p�ȫ�0[�N� ���>��5r8F[Y���2��\������W)���L��{�=�������!�~ň�;��
�wv |rh��!�P�`	CPE8���	-%@Ç�y�B}�9	��M~�̹��t,yBk�hWE#qG2�v�"�mu�j=�g��p�Xa��T�*Bh��	%j�]�y�D��_M;��Kh��ח�D�	p���ԛN.�@�����`��xK#�e��8�	��𑴹���ϧ�*@��zd��#�@���V�qۅX��!n��OAߑ�8�����".).�������gtm~=߽��^�@�p�x�����������O?(��H��.�a��V{g�\댥+�l�#/��}��Ó�Va�����i� D�S���Yd�Vc�*G��r���~����!p$�E萞�G6h�]���0e'!,9���vq［0��	����qǜ[0�Ʊ�x8�9���[O�b���p�����`�T!aG�_���x���"�,S��@-�iYϧ������g �y@��Y�.�*@*c@���@�T�F��R�,���$h�b"C���<2C����D78��@��Q@ -�� h8ˢ!�#��U�J\�D m����]�N����� ��)��̤� �d� M��P����T �"|f�( *P%L�4��Y���)Ca_%��m��wa��$�3�$!���8И�*�@%W�z�Z��2��Ixei�=��@X���ґ��}o�@ZK*�<����㮽�	O&�ܧ����?���nl�ۄ���8�ڋ���/�����/c���(�R���4�Dk��vՄS�r% "��z�	���x�z���I�Q�A���xt�6���/�|I�o�����?��+~��'=v��y0ƚQZ^���ؽ��;�P��ə�0��9Ac�R���,�fn�f��Bof#��������9���}��+�9����}�mf.
귢��Q���Xj����o2�7�W�0ػ�a����	�5&���~=��>�t�u�Й�r�8��v[�0���F��ؙǷ�!e ql��;��`��j LJ�_�m!��H�\��P)�&�F)Yp�* j,�!�D��� j	�ey�KBR]�e,h�E%����G�̉@�$�f��`g��d��a� uL��[OlT<��d�R2�S�ip�� te�V���@|R��+	���>\�A��N|D��3��3߾-A�a�wW��v>���Q�)p)��J��9M�S �9S�Eb:!TΙ�� ���~� |
�^&�N�)��S�d�L�2Y���ХWƀ�!�"8�h��-��k��s��^����S1�1��q��l�t(�w�*7G��8#���nE G0����#�2�25�]�QJ����q/�$�x�&H�.��q���X�(�n�yЏ����P� ��oPw��[���=w����)���T�sX�^	�o�%��,Ʌ'ߛ�����1� �@߿
t
�����PN:-��w�P^oX��Ҵ)Jb�� *���cڸ�>�	A���س�{;��V�����Wn�3Eqx*߀ے�qw���c1� 1:�	�)^���%��T+@*s '60�u׺È��2�Qf����1fgL�q�u1n�3��$�`^��pg����u�.i�Q&'L��`
���u�Q�k�$#n(Fy�toT�݁�~�>������ϱ��X�6l�v&:�WH��3�6G<�<���aH�=F8cf�'����S�46��HrG
��j:���i4�(��3�럣ΰ9E�z�/6G/C��è�߈4�v�`n*W#��	��,y|:Ҵ6�%(��B��=f7�#0��6�aqW���;��;_ܚ�[��J[6:�2ў�\�E0�{'����������q�%�R�ѝ�®r=l����<ߙ��шX� ��g���w �u.
��@עB�V��2�R�-@a�S�z��� ��QDz̃��",�_�{|��&��b?��������݂[�7`Ȓ{0�q>fkq��r�ڄ���1u�C��L\��L�_z7&,�c܎[����H;,��P, t���ģ��X��U,O)�x���Gp�xN<�-��~�?_�"��c�z-2�rq���8��I�٩����	�����S���$���@Wg�+�It�3߷ �x@�|gq|w�{�#Sɂ�O���$D.%~J\�$"*$��R�`u�DE�$`�QBo-P	ǵ�4VY��PS�qc0~�8�3�	���W��2t���������d�V��l��<Z���Ԝ��-�_xd��7�2T��E � �O���,&`� �(/�"x��[D ��[�zS>=�>E�������L{\ T�51HE��k:L��C��k�U�E�F���~ D�uH�i[%�.!r0�3�])
��gTON'�9�O�"�f�.3�}�0�h�(Cѡ
�.��$��X���3N+�����}�8>���}��m�G\b��i�Ǧ"-� I�و��#8PKe�0� !>�A�����w \����@5�=�`��G�`8����%�n*�y��f�;,�{�@����㧃�kB�␑UE ̀�g�,����?���u.��BRf!Rs�P����=(ٲѩfxG�%���eV����Փ-�}�(������~�{� *�� oO�OԢ�X5�v�¼#��mO���V _�{e �'�o=�����P���O��V97��<6�S<���y(�[�x@#��y@}��P��fwڷnp��g�?4� B ���#Rse �1��24�4�LR�!Y�s�@h��,�s�J *�D&�����w�@ȓiX!S�s�*cB%9�H�Re��>�g_)��� ��[���A��N�*c@e�+���>畼�X�D1�O��* Zu�-/t�;����p�CS1n��5n�ϲºuK��7\?�&��(�Q�o�ُ>� ?��d`kG3μ�<>��S���Gx��s��؆���0e��3�/����p�pA`+X|b�H�!��D�:%�yسc Ǐ��_}yiN>��_}��!%+�U5(���憭��PTPZ���\�Vo&dV�����:PRۄ�rD���ڃ3�_��o}�#�Ρ��I�y�.,AYm=ϭG6���8�F`�FG,�sǆ�I�Vnp�&G4Vx�-��Q׳2DGa���-{�<zn��z\�t��qn|�Zl
��X(; ���bw�i]�е%@�� @e[�b�c2�S������B\]���H<���H��
�
d���Hْ���d$�&(^PO��iX.��a��g%�6<+���EPN��$D�,O6�O��ƀ&���2T t��+��~퀥�ϥz{��Q��䉥� ��F��v���_�)~��>B�ң����<�51���� t
;�)M�K :U<�P>���Df	��:/���3�:��')�XL�2b2%K	ݳ��d��Q�*XB�(GJ�LB�d�mO"f�������0��c��;͘�;Swb<	�����ZӠ/�2��0��pj���vX���^\��Ȕ/	�ⱕign�>ї ��%4�7�x�V�����@����MG�^���ɸ�?��JƔ+ �@����;㔐Q%�����1�2%�N��˷-����+@�@ݿq�ǀr���%6�Y���Ы�,c@%WI>��W�{��ǟu�uª1ò�>Ԥ��������9�ŧ�v������z���P��iԽw�<�EXTlƂ�$<Pd�����L���1�5�h<Na?9�F��]I�A�aD�(ayn�^<������s8��8��{8��x�yt��>{�㽸'%VFG��Ĥ�Z��f}o��mŐGL��G��.|��7x���7o���CX�䏩�+1.�#J�1,��sl12�����qU�&X����lW<��%)�p�n`��z���Mf�7�����8�M�������M�E��l�>��Lw쭏���d�l�z�x��q�'|���EP��mF;��8�Xa8>����I���ݞ�#�*����1�;3C�-�m	h�2��)d�-§���_��;0P����3�i��-3�X]���y�9���bE�ކ�A������4r��P����(T/GI4t
��D~���|�>���2�>Ka�O��}+q��2<�o��T�MU�z�E��0��{��c#�)NGn[=�k����e=���ʾ/A�zl���r���8O�ļdO<��'2=0'�O�:�А�Nµ��K����=��=[�g~Ɩ�y"d���!�'{_ۇ�>��}�@�o�m��`��e���O(c@Gl�Ŋ4%�J�=��a�n�CT5�eCҶg(�0@�j�%�5��,�E>�P�7��
5\�} 6z��鴌���%����:��9�jNBð!�j�՘u�up�qB>���S�q���8������Q4��Q 4�-�y�
���>���0\����)��{�pP�]Dм�z�P��K��* ��O�@Z���x@C��-�m��V{y F.@#i��hWG�p�+��xC6�3*��Qn�R9F�L�pR
dJ�mm���?e|�`V\�(�H�@� (�����I�/�d��G�nڝ{ꡯH��uxp͓x�a�=a�f�ڳ���!^{�C�mm�ј�� �r:�*RcB�*a!��s���ƌ� �SE[� a�'�t�j���W���^ZBf<�tHH,Fl\.\��ApqU��`�ե"J�cL6t�tZ�vƲ�������"l�ڎ�����\���b��e <)N~X���`��j�]� �>v'��5��x�I�hܷG�=��_>��Z�>��d>�$�?�]9�۞��/��k�o�f�"�
|*������ T��ʺ%����+��i4!�3��xh����쑡�c�6���hr�˥�(��-eٮ� ����h'_@�,�e�l{L�,7a[G���y�ٝ�(����e�Bd�%8@	�;Ґ�;ɄTA�H��7���� f��2@��
����<d�T TA���+An9
�+QH�@w�a����q���KG+J+��� �d�R��r=��b{-Ɉ$	� ���� Sr�I�/�e
��#� ��d`�9��v�`�{;Q���V�gn����c��5��t�L�;o���+p�-�aƴI�����<�#�]�aî°��`¤	����,�N(*+�ɳ��&;��~�~�9N^8����0g&+����p���7��?,�� h�j$��˂�o/W�f�F{q��!ݿ�]�ݱ���Q�Ԋ�Zq�oF[�.�<te��H/�TdL�Fb6+Cj*�PP^���\�~��z�%�t�����eHM�EEu6��"�� ��,Іhx���W��61��X���!�	W&�U�b��S�d����F��k�b�q�#7���'b��c1�&+<��)x�x����$�f�ܟ}g�2N@�FkX�,���?��p[���ƱQ5������0܋�O�PU+��iX�iX��X��2N��E<��u��j�@rM"+E"�J%,�&A	���+�BT���K�$,3��n�eg���BV����lL���T/l`'��`���hS"�4��\G�e��k��&	�u�J¥x;e��h�A2�:a�����˅g,4�a��h`��i���� ����]�nߌ�rU����-[	�M��A��>��I𔱠�)��E�g��f�@�E͐1��E3�c�1����ј����N�X^G����Im��N�Rk��cZ#��cC�aդ�y�/�;�]��{�q׎$��oƴ�H~>�e\(�qJ��Q4�G��'�޴/	������K��1��	��h���3�;�S��Q+ <���{t�x�)}�m�����xlg\���tx����~§�����O��CY�x����oAP����wh9�.��XH����ɸ��9y���k�/��ߘF��bT_,F����s�L�2\�R S�ˋϋa�~���c� t��(��?H �W	d�A�� -�,א�o�]�6��M��'����kH���+ǯ��>�6�����KcA%b�ev���pLh�ð�#��O����L�����_}������tJ&�/~���e�-������9^��{<���Pp� �(���5���:(���ڞD��A<$d��tBα~���5��=�7���H�R��Ee�ȏ�7���GHC!�p�u�Z\[��u������a�n�If�=׏O~����5>����;��I!��S0��	#�1�0:��yA������S���4��16X����:�燢�ΈmI8B��Ds�o7�ۼÕ!8@�|7��&�J�x�AG��+ð�,UEa\�'����M���iԚ|Л��8G�E�FS�&�H����f�Օ��;t�N�D�L���BѨ�Ae�*�j�����S���=x}o-v�/ْ���,����X\hIƙ-F�&H�ԕ���0�λn	��w#�i>4��!|�Èvy����4ܟ$t�G��|${=�d�y0�?�����x?����en���j<b��mV��u�����Ӈa��6��e���x����?����!μr�}����x绷Q�]�y��07b#����4<��'�\�j-�[Rq�����[��ݏ.��o���#�����j��2<� +�P��
/|�,��U�}� B3t�}���qn�^�)�mӼ�c���p��|l�	�#��7�g@E��P��(h7����*v`8����Z��E��,N����7�fN�2��l��{kcl1�19r(ƍ�¤)��&�U�N��H�E��`����І'��	S]*v�����.���E4�iG��"d� ���B;C����$��W�1[<��U!���7_�LQ��8������yy������"˸OOO�2Q�y4��e��.@�����/DX]8m!m#��Q�cF�8kh+Gu
 R2|�/!M�
�5
����P�h�xD/��h���h���2g��Wf<�[iW��T,ɴ�����v���H�溱G���ПM��F��\:�؁ئ�����s�؆yX��x-��q��Q��;�A���d����#��Q�'4�OO� �z��_�	�j�	q�YPE���=<��7o����G`�Zw��h�և�@-�,�_5bc2������6mpC���ߛ�m};q��˨��FIc#*Z�!�4��d�3c���]�;�����eX�s7,�����c��6�kA������.Ԝ؆�wb�W�Px���'E�zC�����H�Kd߃�!�
o�pۘ�$���|g"�C�E��*���e]޵x�C��e�,���M�i�����x@#Y�G|S"�5��T%F��{ڰ�c���,󀲜���̛K�r���9���OBgP��TPe8�Q�Z��dV�s�C�I�9�Kڙ��}EJƱL�h��tŭ��e�L@cZ��o$�nI@ )@ֿa3oG)��	������/`��?��P�S���2|�U) �y_}p�/� � j&�(s	���Iؑ��� :����:	�4�%3����T8C�$������w�!sW>:_jA��x,r��;�Sn���������G�Fl�_�%K�aŒg����k�c��q�<~,�F���k��UW]��C�b�ر���{�p�b�hThlk�N����_}�W�z}��#��P
GG�z� P�0ut�|A���C�:�>������6�9|/��&�;���*�"�t��s��6#3aL˃�/!�Ϲ�
�:�VZ.��zm]�WG)q��:j6ףzs5�����g�� �����\� P����b��G-l\�y6�~�-� ����Z�҆�?�;������['`Ĭ�wѽp�:�/5�e:��4$�!��HPB>"��"����T2[ S�S淒y�ḑ��������[i �P���aE�DCBƀ�j$�P4bˢa��U�PmFj}*2�Ӑ�ʐT���J����c��%%�P$!T 4� !�~�S�æ����uFhnB��p%��3���t%h�cc�;l��`��,7r�zv�ҹ�e�]cr!|:+Z��X�{:`1T�z."�.�;a~�#�e�3�\�01kST�ڹ/��1�'<��{��[�t�
�+4������:EөA ��M� ����h'�Q�( �{	�* ��iOe_���.� eNQ��˶�w�(c�dN��a!��i<vC�	7��qSO<n���Oĝ��{c1I�>�L�4̇��W���*e��'�Wb��]��kĨ�Pf������Y�����1/0;���	4�wR�o;�K���M�?X��Cu(�Y�w�~��M ���T���&��F/��d ���4��c��B�@��I �A��ø>��@�	�|����	�q��"�9�����"�*�~��E
 ���S e���+�C)b��O�|&�Щ�����q���"����a�j��|�P~~TsF�j ��D�ո�^�����=B�;��g>|'�~�|�a�{�����ڧ��}�����-��|�?����7�nw�t+2#qOvnܬ���X�dݳ��0"���E�x�0���m|������O�_~�O?��h���J��_��-^��<����x���12`���1�6Sk@�15��v���w�����/ǆ�p�^�i�N��Q��\G§=���ᚌ���7��`a�-V�/���3Ȍ�Go}v7�p���~Ǉ�8A#��f���bG���ע*d!c6� ���,9)��#H:9?�G��g���RTG�`7��v�*) �zg~~�����#��	�'
ð?�;�|Ф݄���تw@m�-*�}�-����::�5�K�F?�3��p�.���	�Z��'�n�EC�B7<��MO"-�F�и-C��|��B�є�m�<� ��Dlz!�L��\8��c�-:�p�x/N�ٍ�w�{_��а��v��Љ�4����_��Гg���s���g��7ϣW�{������?Aׁ6ب����|^�'���Tw�59cn�z����|�>{Ͽxg_:�֝M�j�=�7�!�X+s��ی��~�_9��'v"$� ��1��83]��M�K���)�s0���K�K~֙���ph�2Oe��6\�V*�y!�|j��R�"~�r���S�s�`����0������qͰ!>�je<���buFͤ�r�LL��Z<�j<�Pt��>��*���9����'둾3QMqP�F"���_I�����A�Oń�\�#�z�* �R 4�X��U�����7?Ȳ.�*c>y�,e��	:���q�ފ'T T@���-PZ䋰��������B[H�s*�����;b��Y�
l�l��O�~u�^\T�Y�Bv(�
OC`�l�@� �x@�p\֑��EF�vQ�+��T~�$JU����i����sh���<��$8�~�	�/4��hB����|˜V 4&�����ۏ7?��-N_x�����7�h�����
���?�lܱ���*Dǥ(���4��	���'^~�F��Mഅ�#�m�^����	FHh�2����;\�=��Y��_~�-/�v����|e���C��2#4I�<b�a�u����X��7>���މ䊫��Gm�yjp�����A�ۂ��y�?V���k`&W��^.*�m�H����9>��Y��3�G��B��P�3%��"�m���2'�^��r;lK�k5d�
$��T��vF$���vE�&V��!8_��}��챑6��dy.e�.����$!
a;B  ��@�T����j��) ��^�!�;���#��"|����;%�[&��H 5n��&#���W���I	l��f����)U��Y<���qX �BR:	������7�>�}�O�T�xH<�Q�%�A�X�j���:V>+Z|�e �ı�w6��'j�fc���ٸq�4��,�y5&L�Ƃ�����e�xᅓHO6�f�*�[���.��܋i�'b�86hװ!�F���@:b�0�1�'M�]w�[��HOKEgG;^~�E|��gx]��s�0�����d��%4Q��?�A!��������tl߻�~�-���cTo݆����$����	u\�п�0*j��9��aJNGYU-�K+aJH�>ڈƭMx���Q�Ј��d�	�K��INFLb���Ch�Q�XD�����{�"1%���������ǣ�o ��X�~�}�F���u���0�+���Ͱ�SBUCՈmND��l�*�����I*�=N�8)�f\�\	@���	m���&$6��1J��$D���04��R��9	&E������L�)�ot�,���Lò���p���1g�l,�Y�<���Ǝ'.�H�I�jv� uæd�Or�3��Zer�J�#V��Y+�n �9@��(� J=�'��(���F7dX����:<�ͻ����!c�6<���}���h��	���J����H�ES�	��<����A O� tFϥdn�i"���n=���0���(���f��qˎ$� w�J%,�sMZ�����1�E�L1� :����`9�9��������`��5u����(e^P�Zb,����NEYwi1���� :�`|oO,l��+ ��S��_�����@��5�u��܈E4:���+H��*��� z�x:6/�� z�e zu��H�GlS��]�A�+��T��AH:?����x�~�.|�>��7�ç�~�~����)>��J?��������7?� /}�6�_8���J,g�v[^�n�c݉���^���9B�/����Տ���ￆW>z�p�:���M���[x����{��W_�����'?~M���>�;j1�{��Zg{cFeFe:cZ�r�߮�S�����9t���ؘ�Y!k0=�#�0<��|f�� ��������;`m*�Q�r�hף&7�&�l�c�#�7��V�����S�]�h5�Ei�(W-���p��\���[�5l�yp*>2q��P��u!�>t9���-�o�p~�7{r�L =��sUz�EO��P��	�M1N8X�O�6�ٶLl�@m�*c\Н���p�6G+�8\���Z�iN��j#�S��%K���D�4�����չ�+@WM.:���^����lɎFeR8J̡(N��Y�Ҭ(���.|�����ӗ���o�����۟�����D���~���|���"N>w};��}w/�8H=�,�ރ�GvS}�n+Gx�+��x�h�9��xL ���3:;�m��;����*�v��م�]���E* �0j#�[��F{T������WOa�ٽ�.����O�:�G0��q���O u��1a��p,��k�����=Q����� h�.���+��t&hT�U����dp*���Wl�p�}�'�K��v9��=C��VMM�
3�Omz��Z��T���t?�ͧ����Z�|�W#co)��V��ߝOi(BX�d�� 뾥2=�%<V���0	4�~���U@ԯ@`3� �c�A��z �� B�H���h6�Tƀ
��(R����$;n!����0� U�C�h0�N>+��Ŏ���+A�L�NE27$�S�� h �T�PBL$aF�`�6�2F	�����P�J�{�ו	cg:"�$�n2�r��]�M�[#��h�%��S���-D�˝8��I���EBC:և�ᡕs�̦EppB�1IEy��ֈG᭏?��_}���{���� �d��rP�q銵X�f\=$�m$Tj2�6޾����_�M�^�������p���c�Z;��q��/�Z��[������o�I���E���>$g >/	Q������u�R��x�f.�[�0^���?C������F��>�G?;������g[��2ߝ
��tD�����Dv�X��S�O�W��;����� *����w'���T$ Z��?߷xE@C�")#�Bpu8�	��m2�I�jx/b�� ��/�?�`�� ���k��R Կ*�uC����B	�A� �GMYL�Q
�6
�fl�D��E ݕ�̑y% O��?���6j!�)�lt�z%�6W�ʺ,�@s��Ђ�rv��z�x�(��u"� �ؕ��΋ *�1��� �!�(s���z@<#h G�p]2rɜD�.��i	����;rQ�
��GVރ�%�0�y߭X�j-{1qQ��i�F�E���K��`o�����*�
vvv�����ކY�&c���0r���h���1~�}����䢷�gO���'�Λ/������jBQi&�)z� �ܰ�v168~m����Q1�TW���=;w�����%H��AZa1U���^�W�����U�zsv�"L������#8t`?�;{;�Fk� �u����NgoB�V{g'�BPXV���VNDD�0���Iz�otf%�GF6�qn\<��̲9X��q<0�^L�}��7��� $K��}C<��� �7����R�w)��_��� ���5����@�5����!��J�3�	4�ˌ0�WD �1�J�L�IBr5�B����e�QaU T[�į�J4x�i.��k��O���q�����X�n���ov���m���9`���f'�M�t�Jj��ޢx{�����m	BJg�H9c���%7�K���&)�;�p�h|����G��$W��������ڭ��f��!TBp'5iO� �xA����r贄�0U�>E��"��'T T�q�wG��	�Qۢ��-&�F�Ѹy{�?��{�f>M�E��c2m� ��ExMs(�n
&<�^{�=}F%���ɾ��mZ��6��ܶ;	w�Mŵ}�
�Z�Q/s�Dƴk`ݡ��N&uj1�P|_o,6�ͅ��V�n���WN�|���(�w��;���~qG��N ݑp	@�	��}f����@���U�� z��床 z5!S�/(ׯ"�i%|
��9\ U<�������E�����4�����q�����G�����?�k?}�W~z/��]\��M<������+���Y{�E<O`<��˄��p��Q��~���ǽ���=�K�(?����)>���x��q���p�����N��G��zԟ�D�k��|G#��x�@���'����8��s�8�+�~N�u��?�Kw������=���,O�s���q�K	ǌ�՘��a9
|^�E��؄���ͫq]�,��c�\4k�����H�iM��t��|pk�n�`A` ��i�\�\�9hLt��j5�}�����z<|��ŷ��;���;���[�<Ф^�2��(�{}�.xy�	���|��۹o7��.#J�ne���6z+�;=q� z�#;J�h&��冢�������r=���:Z�Õ��ƫx�p=����;6��}�8}dΝ:���=�7/<�מ?���ũ�8��G:����8wt^={ Gw�a�����uk�s��]���;p��^���Y���x������ݏ���o?�7p8|� �ڃ}��w{�6oAnQ�"h{n��������4w<��E�r�+X��9��Ϟ;�o�F7�l/���P t�~#�ͮ((�K?��?<����!�$� �8n�}7�yOpz�|�aԺ;q�����F ]��w�����L�$�i7G�.�=Hih����o���*.�Apf�/���L7�O�l�N��t������ܹ�^�ZM�{k���C8�����1����ϴ�>,��1M�����J��px��«��[B��E�f<���Y"�I	��Kyd{�-S��H����@�8�c �8�� �����@���*��!R��b�͊]|�6�M�j!h4�j��?�C���A�?��G�[�Wuv�|m�7��݃���Ɋ���'�(�]
�PZ�P��"�H��RJ��9c�+�RJ��}{�k���u=L����9�5�;�jre		�����()�r�"���mi�R[c	@�K��p�!Os"#�-BJPL��v$"|W2"�7���f�_چ�/w���&�GCםl �UXh���v��w��{d ʛ�p��U���	=�'QZR��O}�o����+ױc�.� ,���?�?�ܡ�o���k���fd�zx���:z��vt���=���x��~���ox��|q�34��
�/x�� (��.�����q��|�Řn0S�f���t�����c� i[sp�1���]A���(>�	�;�G�El��t��~��s,![��}Ɇ�L�<�r)>d�
�$;�?P{:e�0k�~2t2|2�2��n
x��oh0h{�_ �%3 6i�@u�M�lk��$�������ׁ@ӱ�`��q�F��˜�i�+�	F�˂�T�ꭅ�����T)x��@�����2�sHk��! ��GBK:��r�T��3��`�= �ޞ���"�"d� �)��9	�	��Mq�n��(g��߬�~���de ������鹅;R��G@��ȞR�G�-j����6aX��C����	Jr��d.��ZsC�GAWg5����%p�����ܜ�QZT@��������#<x� {��/�Ȅ��%V/X���1u�L2Uաڽ'T��� eU�7��K��h���,�݆3���x���\�M�7!&�?[�Yb)A�¥Z�s�Ev~j��4� 9;�ɉ�����V�l����
����x���z���l@���~��/����?�_~�O�_�я���K��M�#8,�ƆX�Q��vp�p��$ ^�����a�	HN�F��&�޷���X�b6,��i�'Cs�:�����Zp�w�k�'��BO �']F���������%��m��h3'1�;�����#�, �5QH  �-E,h5����0��0��3�"�5)�'��ya��,Z�\H/� x�1�덀,4��=�0�+������P���G`��B���4����0M��a�6ƚ]i��$m��Ц��0�B�AR j@|#�;_B/;�PN�:���<��6�K��d�^��	
�oêL?L��ĨJ_��싾��B(g�U��J�/Զ�CY��2�<�<��(�n��,�N�>m����䬸*��-�>B��(�m�͞P��Ub:��1�Zi�&i����	B��(��rX��5$C]��l	R�о7�n���Xt��`6Q�C��T��pB$OyZ��Q&�����c�P�ڝ��Ok�{�{>ۏ�_=�@�� �.|����	JR������e���#�v`�w�F�����F�9��]�б�8g��q)|z�S'7��C�wk�F/zf囥�8{f�bX�3*�}�����x���_�I�>��=�����i/D@K&�Z2�(O�Wc\�3�^�o��ׯ����q�ǻ����>��[s1Jb�>����	��%�J޸_޽��?~���;aQ��������1�����z���Bͥ�揇������~y����sv?FG�@3�*�P�l@ԑ:ܤc���B����)�O����Jhę��4��J�C�t�]��5�H��x����%{'�<��:'�g�܁BoN��2	�3���=���V!�y6�]�!�U��ȢcwwZ ��0�[��+�b�xe�����(��j���Y�E��R�G��A��/슳���h�_��:lСi=4���9�m1V�o'����@gm�7�T���f|R��.8��#d���	�y2�hI�;�p~)�ێ?�^ū_��?���O��� ���_㧇�p��%ܸ��<�1>=����`KM*K���P+D��!,�~�����BX�R2���.G��p�����<||�}�1Z�о���QR���H/�4Z��:�1�yf�a&�����h�nD|S6��;��/��ū����/�t�}1�f��/уhŁ2\{t׿��?߁�,	Ƭ���z�0�`���,(�L���$�Mw"�8Y>0���!][�<OD�E ���e�d�ǋ|$�r�!����2�;�0�A����̑1�C Ű�6Gթ�]ۉ�7�b�����E'z�'ÿ� �@�cs�:ɀv��ʅ�י��3��=��C�]	J�a[̙?�C���$�'�!ђ T���§}A+���'!�����/�E��ӥ���\G2�]��O�Gl�����e��VK�ه �G �M�'l�z�W�����^17�oUN4�%%�ܵI��9�ےM0՞���DZE����������h4ڏ_c���L�J�$x
l��F�i_i�p�_��
��\@�R�ƹb���6\��V`�m�Dfƣ�@tϡ}�p?�����S�g.x��~ŏ?=�����OO!����!��M������k��g�\����b�'��q���8���oބ��0x���9�N�p�u�e�5�9�`��*�3]��f`Ȳ1����.�1`�(�D;��X.�v^\���mȢ�U��T�5�%�Λ�S3A=ٰ�t�7o��-�R�$�Y㓓q���@=�ڳԹZ"��|_e��L	H]h�,׉CpK�
�mJx'7 ֩n⇡��Ћ�P�\zv��.���yÉ˱z�������NE���G�A�E���X�N)�{: �@&�f#s� ��H��ɇ��� \G�&N@g��<)lv(� 4{g1����!�%鍹���Nb+���p-=�1��̂ˉ���� �kʼ�/��G�����(ɇn����j0��~�1� /CP�=@1r�@(��u턾ձr�6L�q��><��'dc�ȡ�13BnF
�}�	�7W!(@���~�'O���k;a��6�W���Ƀ������K+k�l��ҹ�0v�����hbT_M��󧎇��)����X����q��)j(ǰ�� ��~p��'������>�pt����3���������tD�����I�I���<����c���y��g�ϧ��5�Q$(��^��wj��߻�c�O�����
�W�� x{K�={�����t����C00^�%�0m�d���5?������* TR, 4a_&�8+$�RG�]�|�8��El�A4�d�EK�	0*<���|�}�_쇨�0�R#�.&�Abq8�K��@�*��T���Dd7d"�������PT{B@������7�g`Q�jAaHw���!t���P*�*�;JC��4�YX�fq6p�����+�Ju�Ͱ:� 4L
��dح
5Ċ`}h���<X
�����.&��-���To��rEb{�<�ߑqw��dj�v�&��n���o�@�v��z��6y	/(��p\�*��y=�OujW,�Ǟ���'{Q����v��W�5�-4�UE��vx]����V4��0tg4��!�*��"�.�g�z(4*5Kh?P&@eo(�B�'f�������/���ET�F:�mAPn�@�z��4T& ՠ����e�,}�	�Gj�x��~�Q (� ����ɼ�q�!���x��X�뇅������2����R ��F�C
����k�
�=���	&;���#һ��Ɉd��X��b��|#��w%���W�J�C10�����4�PN&��O�t.[h���2�[�Xi�ȶKףS+ͧmzl�X�}�r�Q+v�X2���"p�	w_?Ņ{��ԭ�(�� �x�1�zw�����H�0��,J�F�'-8��U|��[��s_>���?}����`�is��ig_捇7q��gh�yn�i�ʾ�A���"V�G�r�I��g�?Z������G��<�}dj���64��mu��=�E����8\w��ؘ&���*�F���d�$=|��n���/Z�,�:l#��8�k�� tOCn�k�o��g;2Ж��e~ؓDS�/@��d�z, ��BN�RcL�v��\�.~0�\�EGb���1�B��r�Z�A��\T�-C���K�1Es�F����Q�
�A��B���*�uh7��;�LuF{���}��@�� �N��`lK�Ş'��u�d�_ݝ����V�#�	�qf+�W��!M�������5<�s�螽|v�X�.��
���]�(�OB|��}��ꋘH[J���&�z"6�$����+�a��XخDh�
KѾs3v�݊��r�d!3��(2N=-��\j\kyn�� ]PS��t��jDէ�����wq���8��ql�Y	�@S�vZ���)�붎�gŻq��g���I�����a"�N�P�9�g7r�c�n6��d�� 5Mr�Y�-ܲ�^��r��q���������e%�����U�����J���6�K�˶;�S�?���Hם+$xW�ó�^��p�j�3�02�mJ�,	:J9ܖk.-A��C��sh��"GX���*��i��V���!�,��IwɞM��N�o''/g���<����F��� ���J��z>� *�tiܞ�ۍ�߷�r2|J���]�N6�g9�Z��\n� ��ܑ=^��PBׁ��ɵ@���b+��d�#���(��Q�t]�?'hhs2�]��%�K@(�al�AO�D"�5J�|�4�}L�iݐ�	��HԎ4d)F�m���q�y'�#��.�O#,�Z���k��NV>v�ˊGB)%y�Y��T�]��q��3�������wx��>�ߺ��������+,�����!�޽��?��+_`ק	�����yZ��ۆ���=L��M+	��/�4����v�.���iD/^1	N���|�;�����q��	Tր�}y�ۑL�����1�At-8_;θ�`��&Ro'���%�z2H��b9+�����8����eo� PN�O�~x�w��4��	)g/�=�����%A�t�ʢ���`�gz�(�Z��nN��CϮ@��
��8����	����)pGTi RK�P�R&�Tj�~��/��3i{	*	@38&=�* �Cp�6Ɖ>��5�6e��x���М�%�����C Zq��=���H�1n[b	:��W���!�Oi�O�8Ā��2���a,�/�
?���c��}�iX�E$�^�0-Ƙ�C!��z(|���T��q=2�2�������qx�:����oܽ��<��$����r���������/��o/�BF��z���7<��=���2N?�mMM��̀��;,tu�a�B,�2�ǌ����0�8,�3�+����a�H�BJbr�㑚L/� O������
�$+Wk�����GNE��"!91q��NAYi.���PZ��];q�����1'�({F�;j��b��΃��v�&.\���G����|�	����ۼµo.���3��T�	:ez���K��3�Y��+Bt+��I�{I/6z)1T24r��BD�?���ȀK ���C�{=@%�@�7�_x���+�C`�?����Ɩ�"�<)��H��H�h)}s22jS��ay!�FX��>	>%���� �@xf�b��<t'������H�P� �
P� ��P���޳�bܺ��o�k}tak�t7��:t$%2����Ǌ��X$��ed�,���K�Ӆ�D�0��ܰ$���8z��~~_�z��Z���)�nU���.����w�4k��AR���jO����-�$�Uk��� �b�����1e��b�|HeR$�Tn��9��%��*66б(�:�}襬Z�C���r�.�g�z���a�
�8�P����1�J�ڛ�Շ�k �ߠ�t�b���h&p��G���F��@0 O�����ۂ�dO\"�P5�����;<��������@e?��P�������Z�u�!�N�!��{��D������>#��������tM�xv&���UBb�$H�����0�Ype�X�\	ϗ�<�����p��W[<����W�B	>���L�#W�����3���wD�8d����g��8�tkT���#q�ѧZq��g���/���=���&r7�{�SR�1��#�=1���i8�>��r=��  ��+���\������ѻ"u�f��@��h�e<�x�(>���(LϱG�4Ch�@����V����ծ�̰��d-fGZ���f\%�}��g\��2��c��!�E�@3�}�7"�㭸��E��ezO��LrC��}������I�L�(z=z����s�1���O�v>BfҢ�Q�掯Nl~<�OZS����*�;��zH���x����^����cD�`�lU�[>�H[��b�.��w�YH�[�L�i�' �r[����i��n+��V�|��*p��7��G-�Y#a��m�����M!Fؗ�g�7��2��X�6Jm)fhN4��,�$�^2�v��`]>ޞ�Ϗ�������x�o+G[]���b��4o����Yh�JGY^4
�"��� [8;������v�M�@_w֯#�)�1�S�YX�a<��Ǵy�0c�@,'(u�6FZN
ʒ�	� 8{X�Җ�;:�1}�\���;'!�gN j�)�ڈْ�;���Σ���ͳ8u���n�u�=f;kcy�1��5[����8{�8>;�G?kAjUƬ��kG`�����I :JƓ�$����)��!�w�v� �V!d<Gз�m ���k��O�d��M����qh�C��?/�pi�� xU�ڇ�Z�\��D���s�\�	���aS�'6��sɸ�! d��q  ���e�%,�,�Z�Y�|�LKPh�� ��Ai?�����;ߖ ��y@y{n�β#�T[!+қe�[�W:'��xr74N�ɑ�nuVKP@�{�u���+�xm�� {��i�!��m��!-Qd������68�#{D���A'j�u��jM��>1�
g�{,����0l����k_&�C��|�(G��ͨ:�-7�b��]��[�ol�3�lC-�X?ˌ���j6Zn���)�%t���.���w�'��C����dde#�0QI���g�7��}����ē�2�`�� 373�`������\�E��;�WOǐ�c�6c0z�S��졘j�VI�(��	�\��g���4]ى�O7!yw&�v���%�휙��C+ٻd���]�ep�K�0.L�@��5Z&�O����6EHa��{W���]�����˓֕�K�7�]�T膀�ķ� tS��	����I�1�I�-t#̄�,��oBp����#\Bi��I��� �I�|
<��lJ��*��t��f���y��X2�t�;� v/w"N@g���/�� �6N���~��\��q��(�঵�Zh��y"n�t�Mە!��ƴ� �n��ON%-���j,C;<gt� ew8g�1�@�>��/}�W�.���C�]�_��4�������Z� �Y��o���C{I��۳��o�q���x�.\� �z��%\��n߾�����/	H�f���_i�w�΅S�bWS#�ҩ�ED�9�l�Z��?KfL��i�h�x̟4zk��� jXoGD�� 6* q�!����=�,a�`EW�禣�$�I�$0��B���		�F`�;�°��'���k���Ǉx��gbPΛ�(�(1a���G���?x��U^�%^�Q���'8��~��[c�����l:����r18<�< !cȷ$ a[b�F/�V~����?*�d蔆�����3�^d�7nw��%T�~��g��K�� j8�����J.��DФ�(��h��(�Oi����D�nJ�@C���I=�ERh g�%�#�.�w�?�������J�zB�/Ah�^P��j�	>{����nP!��>B��=0Xkf��*�0
��u��S]ao��A���w���2z�q��_W@�B���__$$�a�`�V�c��'p��M\z�=
OlÊ4L�r��b/��&}T5HꛤR#���	@U6yA�3�� �J����>X��r�i�@P9W���]	(m���Uh(��l2�*m��X�+J��#��'#��`Ʃ\џS��=7�4|r6� ��-R(�>�*d���zchs�|����Rч�GY�t��x�B�����d��o�`��pX��B�r��ބ3�νɀ�� ��4����~���0�g~�0����;¡�'
��!Gp� ڳ5=X����n�d�X�O�LZ����� ���R��_EJ�)&�h�:zV��,z9�-_���m/Gϫ��F	T	B�U�`$����6ݏ��]y�N|�5R4a~�7F�a;�>����n�Q�C��aEk	��8�I�!�0�o~a ���HG�IpM�����7��d۔����f�k(T٠G�z�؉�Ԫ=��l�1��pj�A�7'q��׸x�k|��m�ڊi��@�+���AľM�������q[��Iv����J�>�'�K����K�Z(��4�O�r\�H�}�߬͗����yf+v���pM$��I�� �*h���!�l"j#�PA|Q�=�C0e�
f.K=h�'��3������T�X�' ��|�٨p^�z��h�'��Y��Uh��4�6X����!XM[���NFY{��FY�!�{���o�Rmd��C��Rx.D��r���8x6%YbK�+jr\P�h��D{�!�=�9�N(M�Ef�3"|L�W]z"����&prX3��0ԟc�y4�]���H j�7t'c��Tho�-푘�`0��@�[:&6+��	I�l�7��|%�m\��K'c��)�j�Ӄ�0���$�\o��~���q��I\�s�?m�U�=f:.��}̥��wRSp��a�<Ռ�G6#�:sMgc��X����vs o4��3�>���(*X�Z'�f�1̉�6!����(�8���p�xJ<Y>7dTs�E��w�J2�J=�Z��Rw8��::Ñ���=�H��r9���\%�3�:
��[��:���ְL# M��9��KCQ����2>�h_������x�H���M�#���Y�,I*�f�(è��<{�Oas�[Μ�Il8��+}ߝ�{�BCwQQ ��� ��M ��^"���>�����>�d��}F�=�ŵ>��gd]��b�$��a���7���}t�P��J6z�w��	�ґp�X�h>�>)EɹZ4�؃�o����6�Bpe$�#���y=�������H!���c��6֘����>L�MaL`j��� 7����.�iW�|CWCy�B����X��f+�@o1f���I˧a��	8w���Aϱ�P�1t�c�����Qr�	�n���`��gP�y�W"�`�'���'�%�g0�?=�d���w�@E�ZC�nF+<���K2tʶa�' *��<�ˏ��E���� �1�AuaHޞ��`P	�Gn�@�1�L$!2Os�}��Ȅ���Nzo;|���@�: 4�<� 4	uy�,�������!�9����\�OP.��+Qx� 0@Ͽ&B��E\MN�O��' M��VJ3�)W h��RT����O���v������eX�A�����^a��#���[i.7��@C�i?ے��;�'+�I/�U6K0r� t���^�1k
������//^��K_�*�&^>'�"�|�+ٛ_�-���XG�ڋ/,�����.���۸u�&?y�g������F�C��__��ӟ���<��;��}�TT���HD�M�0��s0qD?��s�����0�_g;SIܑ���,j����p�pB\Z"����A���+	TS���JP�0j����H�	AaV꫊�g{Nz�/}���_·����Gw���O|�ѳg?��ճ8�����(nGl\ t���`�lL���
�?�� ɧ{T(Adc݇t�m�z���a/(}L��~�$�h٣��螋���x9�m�nz����t���_}|j��W���@D�FV�!�$� 3��������t�I���o�	F�� ��)Ѐ|z�(�����¬s�� ��
}zB^�I���<)�3�v'0��]�!r�&�I�|X-�V�NЍ0��0C�� �ez�.�'�$#�=�%z�
0��X,���<��)��x_�t�G��8��R�0����ћ�XNf���I��JU����h(�N�:	7�:Ӫ��2�6�<��w�.��$����j * ���j	���B0hw���m	��W�#���<gέ�B����^d��g�[�� J�����i��&c��D"R%C��h��% T���{�� �Qj�@���qd��HFȁR䐱�����ڽ@�����E������d ��oϐ�^�uY>X�9SvŢ����P���;�!G��Ypۣ�# �A&{=��PZ� ��a��� J���@�H�-��� �S�Mzn?����Ї�w�g�K�:7��̷��(�3+���� ��{`x�+��9�o���W����^=G�B�L���"o��h}��������Q�ad4�W���_�2(��x�ˏo"ag'�bn.��4hD�w�&d�al���@��
�N�Ze�.�v����t�	,}tಭ'^~���߼x��?ߥc|��C�硃���q�P�Z��ݕ����xvG�9���ۡ���N��@0'�h�n����n��C�a/��.Xo�+�y�Os��R\&X���1����?��žR	�g9aS�.�,�!�y>v,�KP���̘��YF��fV�haɲ�;��W�B����NF�����C��BlvY��%�q]�Z�e���F��J�JV|�G] h�#��c�6���8k�'ڡ:P%���9�i8���'"�`"M�!@o�����t&\�'Ù љ`�a�d��F��r���E�hڞ���d����`�a&Lhhi��&�a���`s	�8s(��k`f����d(����5�+�a�
�欚@�S0s�h�]66���r���9,Wa�Y7oFiO  ]�Y���a(ͧ�\(�'����>��맱��v|r���`��J,7��u-7mDTF����8u�	m;��T�E��1�`2Y�@_�9�e8�s������?4�.���/�F,�����-V��%y�M��E��^�$�k[r��ӜT��ӽʟ�k?8��0p��]�{2�m�DG��Z�	2�]�<`��L�@_�6�6V���L|�)0�)Ɍ� J@�bE�N�Jϫ,9	�'��z7�*k�M^������X�ɼ�6�� P)xZI��>E�[����� /�@'�MUOz7������mK M#�9�C���`��s+wk���9�-��L4Ͽ!B�'C���m ��_]�,��{�	�X�[�Z�;]"9YA.+��l�v���l����"�x>g"jo
���L5��؁�O?ő�'���AԝiDf{.�Ȧ���2��Km{�ڹ��z����q��`��阾j>f�]�i+�c��l&,���Z�1x�Y<�D���9��'���4oF�����F���BtM6�܆ߝ��G�q��l��%�5"��f�*A�,DPGr81Lp]�f�M]��^t-��0LFH�5"y50�rX-��d�0[�S���Dm1�k�*���T����2�^P����r{�,�);3I|\+�1�:f{�4�zQ0  �\;�kKP�Yp9	����ܿ(���uAt�T h��L����H�Ld @d�AɃi J��+	Qۓ�Bw+Ah}bSl
 �I�����(�Mm�CZs�ڊP��L�=t�c4�oEʎ�7I�DP��o��r�P�'T��P�m�D1��q�%'���� m��2�/:��!��a�b-�_�HJH���5�L�����c�������dw2���Ƨ�����/~���������?���ӳ�$:���F�������!޽���?Acm�L6`��~9@�i`�`M��S'��ʥZ07�k#��!,.�-[PFۥ椑R�����$�ӵ�	Bh�?"H~�u�C��3b#$�H�BNF��c��������c˖2�9sׯ_��G�p��U��׌��d��'����߄��X��a�����x2z�R��xu���I )	@��t��#x�G(5���(�R�����ԨBh( ���m1���S�K�(�aE��2x��:$_j\��~�-� tS(�*B^���pĔE ��3�4Q%��H(���_)Р�@�#8�^�y�MG�/�$'���B'�N�N �[�4z��@�� �FR�JîPdivG/M��>�ХOW��S�a��	�i��U:Џ5�i�-��C�2H�@��J��:����!Q�X�D�}��>/2�~��6=ߍ��ad+�� ��>�|ѻC���Rg ��B���ʠY�K'� ��!���D;�T��U!xT~G��qx�; �^O��=6LV���늞�P&�d U�Ed�%)��.PO�]j\EX�J#�mڏB5i������R-���N � ʒ#���B0�N�E�3��a}x}� �@�v�����K����;��$����;�����^�9J�/\�
�����@�y�!Ep��7=@��
E�a�EЩ�=�;��3 eФiM��鎒$0;`��+��_������� ���j�Y�<󼿊�Kz��5��+h7���3,�Y������2w'�4��a|��ϸ��	���'�_�O}f��aT�/�R���Z=��(�����adl#3�����W�#��q��5Ĵ�A+���`�_���+f�%�@%���v�^pC�M����=h�ZC�o� �ˋA��O�G�	^v�"tO���c=�C=�*��P�Y��#��\#Pm8s �c����b� c��1z��=Wah�6�y�&���Unˑ�h��"ܹ�� �c4��9�ۋ$�U�fzo���B��d;�AS�)
�͐�o�@�;�g�Ŋ�3�`#�u��_�)�zaめ�&�M$H� -���R�9(#0����j-T;/�&�%���|���-jף>X[��H��e��K�JqDm��=� �y2 t�x-�#�|\��$�-��#�az�N�;�3VNT)�X3U+&�b�XE,�����5�dJo��3�K�Co��X8��Nĺ���b�l̚6cF��1�0e�x̘?S�ƴ�1�`{&m7e�(L��i��b:�sWL���8�����&v�p�t��=#��{�~;;��1�[��9����ݻ��[�~�e�J`��"��iG�b��6�X�EhY(���.�ۉ�J�-�B�ye8C,g���|(���N�� ���6�V��pNs�$�����"�>�`�g�<k�/�%}���'�P�j�L:�z��&��l��"��Ȱ�5A�}{|�	<��^J�2�6�.��r��v�u)׍�]`�� #�L�$s|��Z�@-S9���d�D[�yX�2�r?�w����e(��tΨ�	�l�P�|Z�@�ma�i	�rwv���� ԇ�ǳQ
�,w��yad{E�HCA���!�!�d(�"���2,�!".C�'l�%h%��+�p�	6B�*��1�4�¿�˳$�%�-�D�\8�.˟� ���h(;��$ �01��D�OF�G�l�ۄ���}�{ z��9|��E�mw"��q���H򇡏����K1u��Y:�N��%31q�<�^<c��c���2Y�%�k��a$J�؅;�73 ��(=X�����p�q�;�w��ԯ�q��)�\nC�ǥ"�o��LD�IE؎x�l��{I�I�}k��V�"���M��m��5�@i�[�&@e�r^��ӯ��y>�j������(/� �7!�t���8�{	 u,r���.<��7����#��)�f�.��-`O� =�v��	�!�BiPn{\���zo���]ِ�Nهr��o� �MGڞ�4�0A��L$�C�7��	B	@#[� ސ����H�(���Ϭ�R �i�$�M# ��Q(ꀦ����M
�U�kE����Hh$Qy'�&Bp��)M<��EIjh�Iļ�83�W ?����.5�<�q� yGK��`���Z8A]�:a��Qؠ�~~>���'hij��ڵ�^�K���K~�=P���G���W��/�O���#�4X��V2VY<��뗢p��׿���x�����=y�ҿG*�6n�A��^��/?;
7C,�13�è����J=�O]�����C0v�0�^�3��">=U�����:�)?���M�+�BTl(�����l_�ԔhT�硢,y��$ьH$�I#AX�RӢ���$����p��0wD��!2�N��X��s�gbФ��;�7�$���@`y��� �p�Zc���#�_:�ǀ�)��ʥT�å�% �$D�n\d��{-<��ɏ� �,�APU0B*BV���0D�Gt�g8"X���k�F������>h�%�O��I��ya��z&:�3�v����	>Y
��BJ�*�ݠ��}z+BM��պCN���6=����P��ű��=M�c��6V��`]�!Vs2"Ni/!�d %���âT̍��sU2�}w7�����}�}�sc08�è�$�T���z�R#�VyA��S�MohX�&�U���[�zUѺ[� ����5��1�D0����z��z߿�!�}"�(����>�B��"��r'1��I�3���Z�6edW���D4IJ[}E���5d$���yb���;r_�+����-�^�n[�ą�P� �IR���5�O/h���:���5���9�Cҫ�_R���*η�(����3��<:^:���_�E�~��'4����0���9�>�CIx?��mO8�wx@��,<�4��[{� PN>Թ5�䏏Z��@XJ�_�	��7�ɀI�D@�����@���0��꽰�>y�3=�]�J�Px@D��U�z��h�C�F_t�W�9�I�s�"��>?2�Q�v�؏7q���$�cE�ƬTw����jKۃ�@ �%�z�r�DF���H���<�!~ų?����_#�������Шq�|�-zV٢G%���;�Ag�j7z�k�#:��B)�G����g���+<~�3���Wn^�U:66Ҽj�0��/�*q&P�^�h2�{���	BO>�
��Ľs@ОQz���.!k!G :&���޶�����x{�@�K��=X�맷b[Y�d{`[�7Z3]P��d�9�4��Y��0@�D	>�������1Wk����l�\,\<�F�Ě��7����H5��<��(���b��(���
۹�p��*�E��X�*���[���u�b/�F�>�(C�� Э�(�ZKǱ���a"<�˼!���:#�l@7�T�i��0{pWh����	�П= ���l�H�h�-3�	0Z2�ړ`Im�r
�-���@k��[���hk������P(�QAO�)P@��}0z�HL�7���D����|*�,���!��7B�fV-ł%�0j�0��O�^�i�1'�Z;��l0�M���_o���+8~��ًM��`���t�K�1��,E\]<�?��o�Ł��H���3-�6��!s0�n!��/F��0�r1� �Lv�U�=�R�����d��лȃ�e�j?�rِ*?8Tp!/�x�y�2��b��9t�`ڒ��@Ʊu�,2aN2"���d %Ù�R���_�'� M2\`��
�,7���� �<���z�V�I4���S�`�l�'|�J��2� 4� 7ͱ>i�=l,ߑ��ɇd	�84W�%틡�4����0I0�q1m�dIˬ`�b	�ts��i����/� J��� ��,��D�NE�����4���HAz�J�z��	L�kD�S_�/�֓ʹM��3�=�l�x��b�0��7y�F§>�lv.�?^��Cx�QD���5'�Ώl� ����w��'��"�7AۣE��z,�'
Q�Y*�ס��f��؁C�O�쫯p��m\a��	׮������1�~q���¦�ۈ7ڰ�H;ZOD�g����8z�>�{�^��_��Wϯ��g�q����7q��m�yF���s8x�S�u���B�d-$6JEG��N^�`N6�J��L�E�n& %�dx�#%���@x���)���[�%�d��?�߲������垴=�ɧ*|��p�]9q\�G�ך��M�d�G�g^(�/̓	@-EBM+j'v�7�vQ[�:���}��n$_�^���PT��f��E΁|�ON"x��ݟ��}��ɻӄv� ���Ն!|K��ό�H#��!+�����|f�f�.D��2d�(A�Bd��t{	����3��5���%��&�&���.��`��nb����^8[����u���c؃	j	�3�M"��%8�C�Щ}�NAv^:�Ӈ��Þ��<ݜ`������55���5<���퍔�X4���ܩS������9�ރ�e��;b�/p��������)�_`_[<�L`���-��	c0�_PQAee�ST�@uM(��BNI��ä�S�gl7oO�eg`��8��y�l��}�{�vه��B$���͢�J<Agj2s�Qװ�voGQ	cd�i���
�w�|��C q���,�`j�3{C���b>�L�AS����%���F�>�F����q!�^bq�1��pͩ���ɖ�w���n$�kĶ8�Ͽ�q�Q�O���^���$�����0ܐ��P �0�E��(%�B`�?g����Ђ��<��x�x"��^ ��K�Gjtv��f/�j(@U]	*�P�P���2A�T�$�V�Eȫ+�����(����!�������֌�B��XE����� ʴ`���]�屮X������4��v�^��Q� G١_�)rB?�:M�27�X���B��5ȨT�p�R��6���1�ʰYM�F��RK�l�7��xXK�VG�	4E��fO���2�lI�D���r�[�ʙq���a i��(j�x?ȷ�&�����R��ŀ� ȕ;B�u�MnP��.�Ip9� �{��pW%U'��'S��aԮ(�k��j�L�����v'����^d���p��Z���b=?�d��X2�����6<|zxM��%�Y�FR?(Op{�N�{�+�����?��zWq=w'�_�:�7.���k���囗��V2�Ȑ�3j{#�HC�m�dt���W¡�=�4�G[�P��@t#����.���Y�'��G~�����>��yع�ב&���T�/�;���������m�6I���}P��7u�uÿji_u���ӹr�OP�e�x/zֹ�|K����Q↱Y�Ȼr7�.�x|�c�\B��2,J����@!CD��~�n	��͑P��ŤT2����I|����R^|�-Zr01�#��Z��*7t!��Ɂ���Jmг؎ �ꅮ�&P2����^8��x�8��wq��U��u9;+�>��Ӝ�e �"���C��a�9��Gx��S�zv�?�E��cCA�ǘ�_a��)r>�^���+0�kO:�X;�χ��<�&ڠ�>���BP�DP���͙v�c��*D�OE��$d8.Fg���EF�$��0kz?L�: V���3Y��3�c�9̛(���~$"֍B��	�ҟ��i(�����(���Bۙ(u��
�(s[�*�U���G}�.�����y:Tͱ��i�J��`6�k&�a�P����0M�+��wÔ�=1}�<�WƢ)j0Y0.k��}�d��NE��D[�C�����Y�E�/� �n�lL��y�' 55m;a�Oq��y��m��H�L���	f,��1�	@g���y�0u��" ]���,Wb��J�ج�z�X�b6F���=�L�a��$�_���Q&����)d��o\��/?ƹ�a���u�lו����t}��BJc�<�_]=���E��̷X��31�t�����%[�����$,�0�c�6�n0���s�|�|Q��}9��\'��r�{wؕzxz���ӊ��|��'��:�"� 2ˁ�ю`�Ax/M�X<n�a����	'2�mɈ6�����"���ٮ"׊@�<�ƉV0$ 7I"(L���L�>ma�lKPhM���|J���D-��o�|�dT�͢}�~m��r~GN���>�`ӈ��0ބ����q�)L�Ma�j�t�d[���̷��y}��m
%`	�4�m���m��dg�PB�1'#���7���j�$p%�g���yR���:4��J#��1�N�
[.� )�=	ɇ�K�рF�R��a�oeO+��-Q��}�8",TZ�J$�!۝=}��?��\�i_�l�FǾ#{�w(IG3�t���X:�N��|v\߅C������q�5$�Ɨ\��u\�7�u�÷xH��#|�i��q_�~_���K���?_���?#���N`ϭ}��u+6_j@��Ut�%����x"��1;	<9�k()��R�����cI��E�i�'����r�Hxx��8�İ)�h,�F��t=H�-d�6FÓ�={��h[���7�&��a��q���tOx_��Ѧ��C���^i�o���L��3@;r��w��y��6��b ��E@Y�3`���{�X��ܷٹ���˭��+�$'�A�{����Y*��+��G���[���`T5�S�gޡ"��G��lf�:�R �F=P)������Ɉn�Cp]8"����#���v h�<��8O�0�=Y�9� ��: ���Fm���(=l2jaog���⾣ jt��'�A��ǹ�Qڑ~ZSz�Φ`�!�]:a���ӣd�q�x��>?u�yH��c� (��DZ|<r��P���M�eh����;���c���x��C<�3��;�)��[���٫�������Ƿ�}k%b���� Ogx�Y�LW+�F'at����}44����^��ٽ������#GBk�<�o�C� ���p��7x��W<��1>���5#� 3,�����$�����������~x�{�C��Mh�ՌʭI���������V-��E31p��9V�v/��YI�Q��
m��!���TJ�qr�$����Q&���4����S�_�F
���H
��Ԩ>���g ��=�$�E�E��,	Cdq��	L9�67�ob +�iP���S����e��U�#���j�$%(�+C� T������LR")j(A^��SU�B�5i~?5�RG�a��#cD~�k�"����H�l0�b3�a�Xn
�`[��1�GE
��>������'�Q}j'�E�c@���A�����*%�B����P,u�R9�&O�V{���հ|��^�Z�*�I��@��@C���p�H �H ���IbO�J�����DYJ�j�}�B1��s0����P&#�k	�fc ������ᐯp�\��	<���x	��j=ћ�s��0���HW%������AF04t[���6�`W�y52�UDh��5z�C(I��S� F��@��C��c�K�%����ԏ+Qr`N]>I��g��v (���b�{�r�I�] �3X� ��Kvh�������>?�����b����P�E�7Jt�:ʮ��F�P��ڃ�S�'��O��ڥ� T� t+'�!�b��n�&���eJ�ް�g�:���P��W�� �wI��D���K�Й���(g��Փ��r�#&�x���i}�_��s�n��wב���}-18���졘`E2X5���L1)�I_��ߟ��ߞ�ܝop�����"�WbV�F�8B���D�+����
{t%�������L���僴+�p��w��q������� �p����u���9�kF���N�XL�DF��O{~Op��}|��E4�AFJ4&���Ft�݀Ŭ��k�%`9�%X�<�ƾ�VLMg#"� %d�7渠2��F���o�3@�Di.�n<!�#�j.j�,�f�oxگ�B��9G��q6.����6�CL+�u� Y=A+�!f�h$��t���(���|��(���2�9�t^��%�p�F��l�[����$�P�徫Q���u�9DŞ��=����\�.���S5zb2��~r�:�f�Q�*Й�6KG�e�x��LF��tD��@��t��LC��TH�{�q
��ؾݱ^[�8p�$}|
/_ý�����s\���؎��*蘮À�}0|� �Z6���c֊i��z:�.��d��=k8����F�1�w�ŚbF�%��`���V����q��M|~�$N^��{k`�-�uXH�:�{5�8/CLM�~r	�o������j{%�;��H��@���k=���J�c)�3�|o>W�Y�1�>�D5� ��Ԡ�P�`rN�<'X2x��4�q�)��a����P?�zt�������j��� PN����CJj�N J iM ��hF���h�`% Ԝ�H�h�@	Z�� �>��<��x��Pi�p��;���uA�{d.ַ&��@�MI&0"'�0�v (g؎X���m��+�D[���N\۔���l(O�8/s�,͊�N �C��G��?K� E��Ɏ��ւ��E�hO ,I�Y�K�@�#�����L�^k<�}	n��8��1tʲ�
 %q�F���Iw�[�Zb9���8 �쇠v:������}��=����i�:���c�(&0.���g�Q{��WZ������0�����(��>������R;�\h�֋-�?߈�ӛQz�e�T��X12d#�p&p��<8	Bo� ��I��F!�� �����lT?�EO�r�'����ۃ ��E�o'{C�Zz zl��C�g�7J�''��d/5{�Y<��ӏ���7�-��7Z�˃��^C�⾸4�C�b���n��hs >@�݄4��g��#�K&[:
��Q���C�',@�ih� ���C��Z�W�P�Rp�QP�G6yBA�@s��h)�!�P)��!4�!t/�$A(�(h�����D6�"�9� �@�`��a��e� 8�ڕ��=E� �R �����m�%H����ȝ\���p�cm&� }W���	8���e/@��`m���:R	�:w�F_DD�굋�y�
�]���Ga��v�����ƥ�gq��yܸzO>ē�=�)��>��\�xW�\��[��ɣ�ۯ��;�ca�|��)�� ��OEL�/�,��lW;K�{�!��^p�s���!V-Z��S�c���I0��u����е���\�nP�.�����P��;U�*q��ܸuW���#Ǐ���ށ~�5�ò�+`mo���T�V���5-u�{b?�w6 &'���0����0o�f.��3�`؜Q"Ø�[`���LDmOF($5Z�z��/��&$���=���i�>By=��} ���[��� ���.	x@��᷅��&���B�@���O@g��S�U�CYE���4�yUE�RS�q��J��S�$�ҋ��CO�^��P�={��9P=��A=�cp��=Gw���^< ���a��
,����`����h��I���ɻ�P�q+�G;�Q�' T��j%���P.r�r�TF��\�@ЧDCP�o�o�	���J�Y����Ш��T�<�����x� ��e�ʵE@UI\�E$+"��2+���I������t���)�]
�ѣ�����g�z�;b��,<W�0�p2p���jd�3`j6��~C0��hX{�p_����^�.ݶ���V�-4��=j]�B������B���m����>b��z���\�&�m�w�?�8C,焖���������KZDk��czsh|~/����8�^[R��ޟ�0��
��H(
�;%�4�6rm�����k{�(=�s[�o�����(�/�̲�4�� �?��u *�����%��s�Jz/�֓�y�I�I9��*����9.>����>}/�/��w�=���qOV�EaL�-&�9@//�;���Op���C����ō_~����og1fg�cD�3���!W愮Ŷ�Rj�����^�nN����W��:_�~���}��s<��	�x�3��@��J2, g���F�n�,+(�C>�H �dG1n�G�{�#���j��A'����b�J�X]���0b5z��c@���eV�L���L��G}���L����+�믍�2���E��dx�O큈2���`}�"1H1!d�������xV����I���Vv���C�j$$ˇ!d�pĮ���#��7	��S�k6�V3Pj;��Q��.�P�U^�QE Z���
�nː�nKQ�Y�+�5�t���0�o/L杻�}�1�/�����5B�(a��>0�
�e#�N� !�cқ� ��c�X�Ӳ��51�og�����Wq�G��Ʒ�r�*.^��OEyY6"�$��X	}]���>��	Bc��=s���iK'b��\�4\��K�~�;
���P��M�8.t#f&Yan�&���}?{x� ��;ɘ?�9��0��"_,�2�� �r\��� ��~׾�g.Gy[�:��0��j�������n>���u&`Y�� 5���U�#\s=�9�{s��7X�8�(ͺ:a�� �;�I�sc���aǴ.{>�i=�lg!�& �/�f�! e��-c$��A�)�{=	<>M���N��' �L�§q��i9�s�п({W��2�+��f)�5�kA�`J2�a�1�������¥�[ g�j��2 e(�a/��� �!s�$ %�8g�e8�qQ��H�)���k���	^8n��DD�HC.��O���+d�1p�׎�0�' ����1>�:�$���,�2�v ���kf�&V�%W�%�oE���(��B�nv\ſQ"]����"����2��q�N�#��B��K�av���#��;^���/�����ߓ��>��3����a�x��D��]�=������?4g�a�tn��/Cg��ӯ�a��Ҵ]3���B@K�J׍=��,�~r]_���&��'�"x�!�dO�/���~�|�ǀ�)P��:Vp	"O�����!t��	@���?����Y^(�`�N�$�6�.p��K��{�}!���E���T!MB� Z�q
�� e(g��X�J���2 M؞���@�R|
 �P�]:�+�b(��]@�Y�~ =&к3[�К���x��M��/�����A-�ts�� -xTXo<�� �4�XJ>��5����@c�
�)~�.��E� �Y3'c��y�]�N��ESC=Ξ�/~y�a����b�����K�͗/���Gq��ܼq���᧧O���/x���.���' �͕���J�_�5˗b�
m�l���-|�|��)���;,�aed��ګ�a�j̚4���о�1�w?�W�0ڵ����P�����ּ����ARr"�46`��]��\��jXQa������!�n\=x��&!�b�P#�H�{����b��72�s��X�O](Bjc�#�^T����V��W�/9)Dr��4����'�� <�m�����:�P���@>}�����#�,�>���/� �0�a@#��^@�EP��B;��] ��m}��1n�x|��	]��^��J=H� O*��@�)O�{���RO�$� u�u�+Ӵ��[	
��9�#���h=2H䇐��@��=�sA�Te�,�Q�31�c=f�[b��5�Dl�p���Ź'7P}r�Ļ`h�>��A����j��d�d((��Z��*�&pT'���E���&�'��A�A�:�=��1W�C��2|� Th�?4��п� �-C��Ebx{�7�0=���A��|��x�~m��de ��y�-������U!Ý��<�ᓽ����@j�е�]	8�3�|���tO�%^O��C�g7���`:��֣��6�8?�!ϾO�NR��J�{��;O� �ѳ�8��d����O�>�����v�N����j;C��/j�@�F[Cу�w�v��m��k���p!�������w���]�y=�n-��K�Ӽ�u���#�_�B����]:��] �A ګYE�z�"W�NsF���F�w��op��C����}s�Zp��5\��h��,
��D�W�����p��K�?p��=�����>���w��i;֕�bR�+qog�#�\�=z��V�C��D�;��v���J�Փx�+��q��W������X�I0�g5E�b`�9T�M�YL�(� ��}���~�'x�g���1�^��A�m��C ��#נs�(����DK�%�a��r,^5��S���ᆨI�Dy�rV"�k!2<��塅��p[�	�e�cD ��&Ȍ5CV�l�a�TL����gb��!<�'����T�b$�V�����X>1ڣ��~<�8$�p�L��Ќd>E�Q�e��P2wm����\	>��d>QU�Co�
��ߚ?D3*`� EL���{wǔ��1w���R�jZOzo�.
W:�5�c�v4<I>W��VL�&�w"#!??�/�Mܘ_��.^8���J���J���0���C���Q}0hl?����Ť��{=�WN���B,^F��9#�{�@$�g �@ߓ����i��ȈǷ|�����G�ɗGQ��ơVX�+ḇ(� ��������_��K�`��6$�'a��ҙ�!V���r64�fCQ"�׎�� CPX���L��і�Nr�Mo�oo����i�E J`i�i��6�Ka�|�z)��*�1�1�u@({99�*���?��e�lx^�������I � ���`�^K�T{��� ��1��%r� �7�*�l��S
���ʒ!����{A��`@�g�X�5J6�e�<j%�`�:�FpD��ʵ7��
�� �h+��V��Ȇ�,n�P�C@# ��goC�L�2x� 4��sop�)�Ÿ�>g��u�Fhp2 �l<�I
�?�ufoe�aKxEy>��v�k��ZF � ��@HZ�@0��0�/"L#wF��0�l��6���|���D�5"h&E�:1{�躑-{�l�}I4���=	�"�kAF �=N��dpp"�6:o�8l���Û%��d��@�3������At�3�o%��-ӵc�j�ɣ��.��0������ǀ �W��!t_�v�Jۊ���,��WKǴ��e�4�ڱ�K �}s�	@�	��wf
�Q`_y�r��� 4��)�p���G���k�\9�{@�;<�����hYM:e( Zt�T (��=\��C��"}�����mI����%�)Ҿ��Y;󑳧���Cqs	Di��4/o_�{t�-8C Zf+��S�o$"�n��F�j=X�l&��z�H��J��.�\b�X�m��r��􂢦T����j��c*�W&�뱳�	���+��OC����_
 e�"H}M� \@���zD�3 }��.�k���J/[��XE �t!'HZ��Z4\ݵz�FpwrADp(��"P]V����c��X�`Ə���}�У'4����йS't�W't���()`�	�ۨ'gG���&�~��ꪑ[����'�!&'	%�H��BdI
��c	�����Fk�>�?����Z���h�oMBܮLQ�)tg|9�T��T����xY4=|/D���C�O�/�J%(��~y���GXa��� �d�4�I�pxe�a��1"nw�!��
�ݡ���ً@�z(�zu{����Ѝ���h�n��r�*�G=�*�z�� 9(�s�<R���>Cjs�Bm�`�6���~�b���fp)MD�����?�����O�ư���i2{��A�ĕ`�@��S������	U%�b e�[��J/���F�QQ?T�M�%%P%Xd U$ U" e)�r�.K� T���� T����J�5�`3������V��f�D� v�t�G�=;Bo 'M��O�Ex-{8L�Z�]UΊ[�%2��Ӈe�R�F�O�k������`��K���x2pr�-�X� qMP%�wo/���ź�D�.CŹf��l��o��o/�R[��Z�k��'(��#��氤��/p�/�=_	�-qX�%�vD�/}��w�B~W(��(6B�9��wk""���JPړ>���T ({9+,�{�?z���ܟT
�2�����?ѿ��۾S����}@ݤӲ0��ڝK�*�B���Q�N�<�_={��?���'����q��7_����=��������焢����JߘG??���n���q��E�}�F��n��N��$_�P�r�b5�h�#�R[� �]#�]��s�p��%\��n?��s�|���-Ƞ�{m�Ӿ&@#��y&�gL�;�*��B�1z�.�[S��N���>�z��?~K�8���G?�ȇ�C��u��V �c���`��Rhn�8��H!��I�@E��%�Hv��T���p��Hӱ�\��k�#�p22�����i�}WCG24��靺h�t�Y:�Ǫ���Y<�+��s�0�/d����H��7�H����79�s�g=���oG�_�<R��r �n>b&�W{(L	n׌�%C{`��)zbR��>=1N�+�����
X1�����S�a�p�������ap\:���N{8��`�L��@d�j�K�uk=�Z���~��k�X�F��N���C1t� �C�^�13�c��t,Z?O ��S�p�T�2��T��b4��� �ע�<1P��!�9��!.�<�ӗ���[8��a��ۊ>�K#�1?P�� �$������@�
c1�|)�N �n6�3�@׸��"ɞe���6��B'��q�pHs�e܋|�wҔ��T
�2��%t�,�>�:��0��d�J I �ɇ�hhB�sH.��rr"�O�Rϵ��+�����\��ᱲ>�tm�	@y�3|�v�*+��J!� �c�����[й�wxAM�̡K�����z�z�0L2�Y��������)����@@y�� �!��j�*�|��O�������?��G�0IC�ba���A��Z8�5�>��z@y:���e앓��o'�w�2(}[����V7�ȇ���	u��B���>�\�1��1�Η��m��-A4L�d��	�I �+a{"�7
���wDмh��%ć�
 ؔ`��D��FJ��2q�0�7e�'���k���^ %P�η��ᓮ� �-����q�a��t?�7F�ztO��-�(��N����C�i[�M!�ж�������5�,��H~�O���p���:��e��N��ha��0z���E��$^y��,�}��õNq�C������[iG�2_�o۳�K��.BTV J6e�S��"\���(<�a�9�;Z��#�o T�%Mٝ���dD�Iq���(iP��V����] �p<y��<�Cps��"k{1rw��G���D#���%ϵ �91�1��.����H�v '�	H9,W��@e	�8���@�a�*����t�rݱ�L�U�S��{+a� M�3cF��!�����W?s�K����^X�,_�iʐ��	��z>߻?�״�gx���ػ���2�v�35���F��e�1iƏ����`Œ��&p�w@j_5?$��u�������.+-5�1o�,��P���
�(u�=�v�bϞ�M�Ǝ�93���޾nHJ�CJv2��rP�V���:$Uf�3�^��H��Fy�&xE�c��i�3ut}ML�LtK�� l{�wċ_�87�,׏)�3���#C�H&u4Ox@�s<o�O3o'�C/Vz�}K@K���� ЀB"��(QE�%�-�DDQ�HN�˂8����<Ǖd�
 ��en)��`$:�"h�L�
A�W�f��@���r]i��H]���C�PPyz���Ba�*��"�|U��X�O$#`��,����a��R,2âH'L�0�F��֯N�ҳ;����z&����tKh��@��j�NP/v�A@��^�.<�*��7{C��] hP��z��*<�^Eӛ}	T��Ib �-�	徢��i�T�y����[�����n�R{�-
���8��T�֕�����n�\`���o�|r(.O���j�:�ծ@I��Ĳ��>h_��̹\;����fW� 8�I�E���cO�B�xICy|0����>V�G3��E��i��3{p��Wx����_��/����]Z�W�V������(�ёС� >g�~E����#l=�N�XM��t��F���P���Ph	���� �h@�mRu'��k&K@��>����s#ã���	�tLrb!�P)P�N��A��B��>�����Do��̱:رx��M#�NlK�x�������Y/O�:ջ
h|W�o3\��w�%P�:֣a�zo�	�J�)<������P �g�bD�
����?��˧�J�y��-�y�~����7~z�;��Ɠ{���>n����^��+�p����}U��a\�ѱ��oK�;jKN"���\��9co�1:�.ƈPT\<���=(~~�o���էߠ�p��b��*%��g	�R+t+2��k�.���K�M��y	��9��1���#�|�/�ބ��4h�-@o���]�nk�%|� б�Xc�u���h�8q�����2��a�R��"$9�D��D��犾�\����kM[O���xX�MŚc0p}�v���)X�f�O상#�1�W������`3g�f���P�i�F̚��_?��F#���x��Ld��F��L�,����j!�z.�,g!�d"t�"`����ÉjX3F	�G*`�9Lԓ@��}{bf��X0PK�*��@g�:�g��ż~���vK�r� ������z�:揖�̑��ўwGK�b��%X�pVi/ņ�˰a�,]4�gM��)c0|�`9 �G�����1d� ��23M�k1���b����=gAz?��E�Ѯ�1;�3��1��r��>b[rp�����8��n\�}{���x��>�Z��NXD z��iܸu�i���<hYi��	h>���F�LNwz��E�FT�Y6�	7�~�%L�� )F�<x�o�Q��2DO����S'�� *��Z�e�)�@	@Y����p\����[���P^�K��@e����bKb��S\&�3�r�!�;P�p*<���e���]�d����~��&t~��Q���h]in������7���!�m�B�:(�' �"�D@yJ2X�\��qV\�M� ���'JNٳ&BE�dN�?�� ��|F9��S������m\����l@ך �p"�q?EN��Kv����	t	@%�>��fdcxo$��o���s&[C�J�L�,�|��G�&�	|[i�=~�	��ӵi'@�F"���~��bH�����|�#�C������md{rX0��7t;��F�M6*��}@��6�2��uמ�����#<VB׍�oHc,�8�=��WAut}��B��zu��t��.�hY�|�q�3'"�d��瓁ss(	hy�(���.\'��[$�~�.��{��'WT8	��s+� �E��,Oؤ8O�k�ϟ!�E,�bO��x�������-.<��o7\�*	@BAG\�r�ۢ���ǅ_�#�(#Ah6ChG(.'#bh8��A_]���L����P[� P��v (��$D�{ˑ��D hf+�k+B��[�٣�o T�4� }[!�"�ɉ�3����b��� ʰ"�D��ٙ$BpC*���j14Ǫ��Jh �����Q1u�X4l�$[�v�Ր��?�+�|g){>_�$c������m��;�_VsP:�۰������}|��'h�Ҁ��lDG�����^���N��iӱh����`��X�x)��H ���j���9?���(.*@~^�|���d1fL��Ic�`p�>P��];u�"VoME�?Z������i�(k�B���ԗ!8#!^pp����vX��pz�"Ӛ����ڝ�Pj�t�ހ� �`1-���{J<nw��P�ߜ�M�=�����8�% ��_��HT(J�$T�"ySR6'!�!q�1o T���CuY<���4o�e�
 �p:�u=;`~��r�I�r�ѵWw�L�� h�@{���O��0�T��2\�U�6� t�,���3��k6�: ��a��d���x��-|���]8J� ����L�/r�Z>�� �� �BE�P�O�B(�:�/���l�&��F_R�
/hp�P�� P��!���J�� M�OU�zҸ �Mr��"�I���ч�=�è�������%����=+9L��	*9���v/��N�*pB"L{A@嫜ѓg��n�C���h��>������T���u\���uP x�'a(e��(�p��~S�|��>H��
Pq������/�����xI�"�,',�k{~�P������S
�|<�#�zr_���Oq�S�>����-h�ĸ���C ��;�zKjŖ P	�z�G�k�]��K)�� i���g�F��S
�>�R �A�̣( ��q\�e�����J�i��i�X}@���+���2��y���2X�Mu<�>�Ҽw��%@�/`)տ��������V뉞5<�@ώ�,��,D��;��.=s7~�_�p��=�͟��wq��{�ꧻ8��[��s�n\�W>é��q��	��8ꎷл5Ȉ�j�!�n4���:B�ږZ�;�]!�n	�#�T�!ao=N��
?��y�_�ѫ����6���[�\܅�IN��
�3,ћ�mK�ѽ�=J-ѫ�]�ͥ �v�	@���{D﫛d<eA�|4<WA>x����Ga��+lF�oĲ��X���c��$xŇ�,�%��(�A^�J���G4�f��(x� `��
�J0��{�Ѱ3�����'���a]0��r���8w$�VG��=1w�"����0�ڏ t �G��H����&ů��i�4��t�iH3��,��B�,� �t:b�'"��7��f����0��&k`�8���9��1w�<�H��(
 ]1Vk&�Bw�fh�piv���u3zcՌ>XD0;c�f�c�U��hCc�X��KW`邅�?k:�M�q��a�A1z(���!#b���4�/��O >g���eӄ'tΒ��c1b�@�N���#0�a1&�l��(cL%��I�$����	@���m��bs[����sƲ@�Ϡ���Z�X��׎���8rjJ����f����W �! ��� j���K�5ņ`��ӃY
��ÿ:L���s?a���᷺I�>uY4.�e e�@e�PYP��>�����ԋ1��(6��J)���$9I/3�1�A({8M	.6eQ�$��zTy_�����&A�;�iM�� ʞPP��k��j�h�4s�������ۢ|���''#�eĕzB2�����@9A�*Ck4��R�J@H����O���<��<��S��c�y�<�MHnK��NYK�d��˄8o���:RIhNN��G��z6p�n �g ��������z����X��=��^�t�[�H��j
�ws�Z���F`�Fׂ��wk$)�DpI�-� 4�/ٞ,���G6(��X�!��Aܥ� ��s��ht���+ON�$J�l�a��P���o{@�24�� N��A�m$�!H��% ��b��|F
@� �;�a��B�^O�� ��H��9��q�"ȯ��(�s���@�lOG|S*�kSZ� IQ��u���}�;2=DP��:�:�{|ztz�P��\�O��!��#�g ��Z$͂�I��E?� ��O �yA�h��4ĵq�h�IG5��fHK�p"�M���[�P������ ���)[���Z(������m}@�'������d���}CP�vxA�BI�%cP�R<?�X>Z���qj��}���@�a�a���3v�}���o�R{�_���w������
����|��4Ox:;����7zk����C ʐK�O�>�7__�㸊??�m�*2Xоx��޸�3�Oc����.�DZl"�]`ed+C�Z���fb��X�h	lM̑��3'N�����Gx�ۯx��7���G����57�u�T#" 6&��!��]:�oo%�k(�� M����9S��h�}\�����&��I�Dbi:���Qgp)�$l�Dځ����>���鞰wS�Tx3�@e?0�d1lzm���y[�NlO���s�-˿�����"	QlybˢS��L$n�g�`������=��'4 [�8�z�5�c�u@��}�o���M���T��b_�T��`�V��0��V��D���М��ak�`�����s�;E9a��K�H��ٽ+���[l�x�y��G��%���@����^P�*	@9;�RGb"M��Y�.��}>5	>���^��FR���*=�H�lr�PUN�jOQO����V�eH��f��cXs8F�D`$i}$���`� *�6]K�Х�ݪ\	6ѵ@f��:'J�P�N��Bd�� T~�+�W8O'�)��f0A*��*lr�0�v�uEO2�{�
B�:��������`�����XO��Oʱ�B�_؍�W��νKx��-���}j3?��kQi�����G ���}؏�M��_p��i�n+�^u8�Їw�(�k�Ǝ8h{T[����I�س��[|ѵ�]Z	2	<��)�O)x��� � F4�HyZ�<d��M��b�;�헇>�|ڦօ��W�Ѽ� �e )�V�T�w�' ڹ��2V���nrGW3�~��L.�Z$!���\}� g�������§�.!wG-��5���64];��_~�/_�÷����/���Ϸ���Nzg�a��.��q<����:h�������}�=��lbA�=���)y��3|{�:n<���I��%���
�~s��o�IE�^��%NP*�E�lSt�2y���1���(�r�����-2�r�T�M�A��%t5>]��!+1 x-��b��j��0Z��А �g5�	���u��I���8�VSh8n+�f�̦+�p:A��A�7�K�0��F��]�o��VOŢu�1x|��cwǜ1*X3�@-f��`x/ɒ!X<�K ��%a�X$�q%�N@�q��T��LG
�h��d�l�H��c�d8���q�%�%�8�Vd.']6F�F)A{�
�G�b�heh�S�j��u��Z=Iڤ���1�f�QÔQX�`&,͌�a�:=�t7@g����OŨ��0``_���6N��}�w��# tԔᘪ53	>g-���F��G�1`��_�ђ������e���`|��n�xǾ8�]oCVM&�c�eX8�,ߵX�ћbq��8��^;�����Vc��T���@�隱T+@&��Ѝ��N���I���Gq6�˂`��@ J�o!Bo���� T?�B��$�d�4H�!���/((���aD0igN�N�����g���<�!�Ci�����+n�����W^Tڞ=��2,�}�O�oh�.'#�0`p\���0ܘ�Џӣ�2�~��K݄4z/���W��H
�<$x���VI�Ȇb8�[N���>�����[�
$m%�l"�$7t�4y:�l� b�z�'�˟*�O���� ���	C�O��]+}�+9S/gl底��t�����u��' ��s��ɽ� ������ݭ�������ػ��8��8�sX-%-���#��0Wp��X�q�>y( �����4�0�A�G-�s�澴�U܇�=��d`�#�$�i�"�LD��B�R�余�ۙ" 4���}݃��x��{�}���0��>���4��&�}�M��\*�[
������=�Ho�E��L�W$
 u˓�)���n��({@����H8$�O7�L�����]	p�i�A�~dWK�$͂��7G�a�$Dz{(���� KF�I���t��������J=�,�D2�����	��H-�@sۋQ�I�HB��4����h��B����v����De^Јvz�聏ߝ�l:gz��9(}�>�28r ���qSGc̄��]��z�"Z�ϥW�ʰ{�6l��Afr2�rr������w�~�g?=ŋ������d��q���0�g]�z��Q�����p��`wK޾�_� �J@ʙ,�!K�_^��//�Ա���)|q�4�� 3)A!�!���]ؘY ��UU���m<��V��o�˜p�ן����c��Ŝi�1a�P���~H �Q't���?@��0c�,X�����~H�Z�Q��MAڎ<���E��d���K�M�T���x|x���Ey]���{K�;
%� T�ƹ���rPYP�h(��e��?ĔE�0\p���!TxD9� ����d�&{JT�>�c���~�"	�=�*ʰ�S��p%(�A�6� t
��5\2c�'b��,1��$G,�v�DW}X�F���~��yg�]E��C��	�� �$s�β�F�@U��T
�ƞ�RPW&�$�T#C���:��|Vz
�T� ���b���P�N�V�i%T�<2������!� �D����H�n�`ګ��K�hg�N�|2<2hr-O�x���b�(�eh�R;��˸\I�y.�"_�"
��ո�[�zаA�U����"@�'(Q$�\���%�7�C��S��a�+��KP��V���=��7O���g����x�A�?!����@�?���wj���xFz�����Y��h,���/C�á�-������P�n�b�/䚼Уً`�][|Ѕ@�s+�۔���t�' *Bf;���yb~Ǵ2E?�/&��� *��ћ�vl#�X�������,�ѿ�Y��濪�]�d��~D�&��ڮ3��0]����Og���«G��/����+���y|r��4b}��"�$�޻K���2��!���!��9���×N �,b]0'Ξ��a%n�O��ߡ5�PK�ƨ��1P�9}�^����~|�����;�����v�W~���]$�)	�1:�"L�c�Ds��Y�O�z�@9����0.�y�b���ׇ�P�-����,G��U��
�B��a�r��ic��*,v[��'b��>X�=.��@`��.�b;��S@��7�+��F��f��`�*��-�;��&�PV����ՠҿ&���Ƌ1q�H# :�'F솅4�3} �����Ap&x�X8��!`Q?�-���#�z�׏E+��qbu�#z�XD�#�|$$���s�`8k�՜~��7��c�$U�����+Ʃa�(,��e4����t<�go�OML��ɣ51}�lذ��X͹V�Ŋ�:X�t�q(���9c*���>�5�����}�i\��Ԡ�WT�xo��<����9c1v�0L7�G��7�����0�q	F���_/ t��2������8w�s���1�ѽ�>��Q��I�i���FX����(n�ŧ���GQ�X�%�k�I�Y� �.�M :�G&)n�n���|-���*o]8ex"�)�%dN@����v+��)�}�n�7�!A�i:'"rɈ@Y�\����:�����g�=�v9���3ن�q2!ږ��Cn:F�bͅJ������4�O�YP��}�r�n�4	�����h"��r"Ѝ4ܘb��3pr��}�"7t;A"({@y�# �����p�O�#�&)4�N�G�!S@hC�@���g`��Ҽ��D�"����}OD�U�'!�b8�q.򗾞��c�] u��iS^ε,	��i�d��	�Jh?�P���!�'"@Փ�ӽ�`�K�x�7C8�T��,/�W�i�$i�/]��2���2o��OP-�@ܯ���f�Pe��{��ǵ&�4�Fb���+���>���AFD�2��2iw:�>.F.1ZdK�����tL��IHؓ�R8��t�����K��ʻ��`�u��v����Q�W�-pC�n)��4� �:EQ".{?���`�&͂�Z�۱��G��� O�?���M�t/݋=��@)����D΁)F�N>��\|�IB�V=�wCp�Z�ބ�
�$�8C���t>Hk��h_-yH�{@�|ڂ�?_ �%�t�b�!�@9	�b��Ӝ�`D0oC(���,�)��0j`E�K�5	�WL�d4�jbИ�6a�M�YZӱa�ZTU��ֵk�**F��?�SR�u�f�UV"/=��,*BY^>�

PQV�����ގ3�O�F/	Fȱ*�����m/ʵ����� yitM����`O{��9 ���y�8}�0޸	�F� �ο�ϟ����s�N�8��{��ȑ#8v�8ζ�&||����%n~{�ֽ'<��c��k�e%����:�1u�H죎^ݺ��N�����г{w(*�C�?}������EpvFX~$�2����W�=����Hv�@��I�;j���w% ��)�`�d���?Cp���~Ը%��Be�&e ȓ�?��td�!(��eKh
 ��~r�mH^� R��r"�DW8�x�9�#��.��BOy:�@�)�*�@w��"�R2�k���"��
ꓔ�1U	��kbĚ�j1�=��,D��l� �S']�e�`˹C8��k��[?�M+_���bd�%�f[C5����P͓��:B��LRȳ�{W{u@(���$���C��H�ĞO|�ǒCmyZ���C��;��,e�F��O���%�C1|k(�q�|���Ma"��g)Ad�3�T���rGt# �h�\���a�/ૺ��o��w�Jww� qww������Apw�@]�����-uw9����ٔr�y��|����r�3ךK��9�c�)��"P��1
�*�)"�̀�}Ű9_ �é0 ���s�Q t̞(��°���r����K0o��� �f�JG�G@���HE�I~�hľ'���O��k����O�ϯ@������z��?�<	����q����Adt�ë� ��@�ρ���+��Q�#���;���}��D�:��G	IG�=F��L��y>��=�����[`�� ��%�� �ڠ}�@�?�]$�(�+�⺲/��ރ���� �N�T`�����?С|�@+�#����U�"��H�UE���3x�@�.���7_B��GД����p+%TV�af}<��x�(^��C|��x����G7��{װ������0��-�{��aX�j�tW�_�O��?��g��O�㑷�D��^��ơ�!/}�"^��Md��ar�;,B�A�o)��.���y��uA���Zh&����<��M|F� }�w���:^�訴���
���cP��KX��e�����b�c�^�o7dE,EN��E.FN�\${�"n�=��� l�9��w�!<f�����^�m����}2Vop!p����h�\�K�a�K����8��b���>ϩ�i��9�������� ��,5G�rK���79�t�$��G�z{P�OQ�[��YK�����&"l��f��c�!T���XᤉeNژgOu��",���|�����1���`>nN�X�`
�l_� olضk7oŪ���x�2,Z8��L���.pt����5LLalb Cc��kC�X&Vp�j�i���:{�	��L`jKX�b��n��\�xAg�z`f�:U��k���K�⣧�܍���b?6&m���J��� �2<�|�o�x/\u{j�8x5��̈́���[ :a������cCA �f�`i�L�[�Y�Kx�hh����K��@Ua����?}�
��Э�Ī e<P�|���JP�����K������E^J�M����  �q@�,�(�J� ��ܭ�^
�J���xB%<W<��*�g����ԗ�ʀ맄��T��NU�T����ǩ��fʗ�y��<�*C��T�S����W���TIBԟ���%���v+�m嬓��Q���c��8TB��A�2�'m�����,C�	��ɪ[ ��/W�PE{U��R�,�@�x;Չ�$�V��H ���pQo����
	��\G`�R�2M�P	Ǎ;���C�H��p(�J�2�zY'rO�ҧT�#Ἁ�%#�H��K�c�<yNI�dB���MU��I$%E UK��*!�ք<Ż��T�1+� T����j��k������*�E*��k��s�e�>��/�E'�Pq���s�'Ky|^����o�8A`���X�,�x-e\W�x�N�R�+ Zy�eG�^۱�ŊT�	��0,��iKV��ٙ���n�'!S�����zyox/����@U!��Tq���7a��u�aX��r(����T�G�\�W2��0,�r1r@k T��#lJHn���TyBU4]}�	��	�'w��A�X��}��
��(D/ڎ���2�%<�R(o���s$�/G6�S�r���+ �, " sd%gJ����55�p>Z��F��]��mi���6L&����nvp�挹�硦��?u�E%�
CFR:
�
PUZ��JB{]3v��c_��g�v�������Eyi�����K�?�O���,᳴ )GP$����6���&	�h0����p��Y�6�xe�(�JEfB2⣑���@��#/9�:��}��ɧ����oJ���ۯ�Ⓩ>����O|��W����x��|��w�叟�˟?�_�|��>��o����$$F�jG
2Ӱp�,����z�9l�,agm�1��``n�M>[�_���W�:>č[��mK�U��ƭ�� ���GW��7J=�7�^
�JܲK5
���T����/�H��B	���	��Lhz{:���Ԋ�@_�d�hZcrڲ�ב�2��Lh��.��/lm�J��m"�ca=�F�:B�N�F.	�����T�z�ё�%`:�%t��xh�jA�R�l�C�AZ.ZЙJa�6L��a�f����uXU��������5�����O���?��߾��W/��K���;��[�͆@h��VAT��8���Ԅ�Ph��������W�}
�j�T�n{	g�R�'I���&�v
	��	u^Q�^�k�/Gs`z0G�aEY$���n�R��:�S2o
�FbpW(F�b��p��	Ǆ�hB�xQӠ ��'0��@����FF�����L<�KHM��>B3AU����D �G��F`$t���T�S�i���o#�j��a�蛀�PB����fWI#v������~\|���
���E|���U���;,�HR���^�G���oR�w����?I��7~aD��P|�%���?����FbK!<����σ3����
`p��gC�dt��A����X��H�#�$EP%T6I��a�\G t� (KB�yB�"U���"�CI8��X���G�(Y�@�^�]��T������Ӫ�S��sK
��s�>
�Xީ��{	����H�L��Z|���H%�НR�S��]C�L4lo,F��'��)�k,��9�n
�uUʞ=��#���|����vcqA8�������=�H�2?��x�����z�~��~�>��[��g��/���K�!�����H���7ͪ,�w���������lw^z�<��+x��U~�(rk�PӴϼ�^��|���^�@��ݨ~�8R�wc~m"r���-F5��Q 4�}'a��ミ>������*�y͇A��L_���+0(c)�,���0�]��Q�1�{*����4��������Ԡy�'���G�vD��B8�	]A-�B�2[�,���Fؼ�����^3��=s��@�r8����i.۬馰��=�!�0�y�^ᤋ��z���:���ș��'�&H���ѕ6�Ya��n�jEyklQ@ (���d,2C��q��� |zO��W-��4+5��Q�𩍅����9v��i?Sm	��Z�3k���vX�v�yn���vl�܎���X�b%�͟���f@g`� ��-��,`ec3K����� F�0��S#L�F�[8S��30��Φ0�i	�S`G�O^�I�1-����=��_��7?~W�>���w#�,CWb6�紤5p�]g�����K}x��kx��GQ�V��A+��36A�aH �aX4�OƸ�����=�.����AK1?t<���Ocw>B����`�WB+����F���&���2�g9�˷���&Ar�E�C��Px�� �O��'�y7x`�Q��@�W�Н1���Ւ�V�+�D����2���x�* * *^Qu6\Y�xNy,�K�'T<�w�?�؛༝`��`�A��(��g%���@Z��i�2������	r�T�}��x� D�8��"��4��R�tDv')	h�	B����X����.UI�X д��P	�݁t�h*�ER�uDBp˕\	�Uy;��p&0� ����y���@'�CէS<����8�$,�@DS���D�J=Z��Q@���ʣ���}V`6CɊM; f�G���z��OCT��+��J��2&*�S�s�H��}$|
�R�Z3]7  ��IDAT�J3]~�x=����L��J�$��JH+AP�_s;�@�N�� hT�yC��*��;V�eѲ����������)a��<�4�o2�a&�sA8��QH��q�%]x�I���9$2E
�:E�ܗH��]��9�'	1݉��D��^U��A��
��G��j��y�nLQBpCjb\�d� ��HQ2�
p�u��6ű.��pۛ�D����t�i~G*���tO��`�H���p�A���{�^Q-U}_U��K��P���;�ڟ��CŨ:����<���R��Zu��ԪS,Ov�t����x���8��)�.CɱR���T T5K�"T��nR<a�j/� �f��=Y���*�@���&����b1���|�)�l1�͑��)��om�;7n���q1���؁��#�
1	��I*BvqJ�:�UT���D�y#8 �щ(�+�����-u;q��|��4�T�0������I�+�*����w���ģO��G��?N=��>�K����������4Tg�����-8{�8�{�	|����W��J���I�U\�%������	?��~��;|�ݧ���<Ё��Jn�u�G_W+����Ͽ���}�;l��<�C���� �U���-��@j��KR���%(<M=�Ʉ���&��=M<׬��x%a��S���$!��*�[$�s���%����$�AO�"�w�#�=�-��l�EP-���p�8F�1HmIGf{62;(�ٝ�J�>)s��D
15q*	AHe$�J�`=� :� :vF��x>o�'aS<��L T�t��3j4ƌ�̏���c�eA�р��8L�4ZS�4T����r�=\�gaN�r,Kߌ� Q@��e���F�%u�=f��!�xL�.\��m��2�w��2j�r���!�;M5B���QK0��á���!���D2d��C0%�J5@%���i���hh�IT rB{ƷEb$v��8e|PU	�5ޝ����`|8���|��Z��<!V�7�;C0�- �tcH7���`����h�n"���@��vo*t��x�'�ݛL8͂ݽi��We���e�	��G��V���`�����D+IWd���-��q��I����'
��	0?��ÙX��/�B��ā���WO�ܣ��W��=U�
��ǣ�D�S��\�w��EW^�;��;�]*�UE$����M�G�y%C/�3�0���o3������>��}�z���TcsG�ͅ���T�$�Й,��d|�1��0�X*F0G&�I��%�Qk!t(�RƸTƹ�c�v�/ ��5�*�A���%�H�S�R ��'��@*�D���#�*�l{�����K֗�8=hO8A3���NqݻyKE�yI	���!|�"xJ&�|w�D��=�1x5ka]����)�$��~~�G�0=; ��ba(	���A����p�5�`	��U8|�|�o�����/>��?��w��ü�D8&���!|ȧ�[��>ŵ7_���^�37_�7^��?�'=��o��d���G����3�#�1�_�g�j�L��=`Z���e����s?�M��7�� �}�*;�0�w1�S6`d�2I[�!��1"e)�$,�^�B�D/�K��m���%Ƙ9G~[��<����1[����Q+��x"|�O��|sx-��7A�w��7OA��g�Ll�����uӆ��(L���E֘���S&��d$��c���u3�'lr�m�4��	�	�w�D�d�M�G�\$/4G�b�,���H���"s�����"~�	�g `�<]d�<����kb�$,弄��a�f;��Zp������,X�����&|nݬ�����+C�-^0K����s0g�TLvv�$U�!cL�6���!�Eֆ0s��)�yfN��LG��=l���d�%gZ@���m�m�j8f��S�X�NŪ�M���%|��kx��c�}�E�XEN[����0-e5�ǭ�_�?�߇W�~���DIk�/��֩�����0�����0=a=�+R=�,q慯²���*B|k::3	}a�HhE0��ckY�KE���X�M�~ʼj�K�����$4V8����peگ2��,����6�y 	zܗl�]����7�����k�PM�P+ۊ�o����
�JPO°wU0�W��{7��'�6�|$�x��n�����Rꍭ2.h�/�+|���^M�
p��VN?Y�4�g�1	'%�#|�M%0�?��Yf���=���N.!P
`����C)s%�aG���$x�ޒ���f��d�%�rY�ABفB�c�t��(e��D���
n)�P�����47�X����SC�x@	o�\W��O����d^Y��@�xQ�h/���T�S���(p�x O�3�JL��Jxp�xjo������*a���,^	)�c� �J>£H��L?R�(U ��/�Ɓ�ⅎ�~�TA:��*��ڲ��kEʴ@3���T� �� *��y'�y�ʠ�#�Wi++ó�w��g)�4��e�P9'*�����t' �6_!4�lWq�e��Py�E�k�D Mh�@bk&"��nJBB��NB&m���4$�r�>�0�@0�D��Y��L�h~O&�;
н�	�J�� 4����?����g�.7� ���:�g*/�Pt���s��'���&p���j��[��)�;�|W �;0K��Qp�;�����r7 o���� ��$"��{��v��O�#�:\�/���1l����b�IS\�4}
jv5��~DW�l����T�K\>"	�AQ|`s��]ք��6����'
7���7���8x�*+���!�ط{^z�E|�%M�����L���B�/��SLJZ���*�_�������ҹ�x���x八�x�Zv֣0'Yh��Ņ�'�����/>�?�ĝ}��J�ݿ�?���S��_~�������GQAB��^l��cÚ�
Ƈ��������V6|�~�Z<��J������(k-B�v�^nS��"�g��(>[~W ���;%�4�ۖ\�T���RA(_P���+ �ԕ�T>���HjMFtcB룔�Ʒ,����Bbc
��b	hf�e*�ΗL T 4�9U��P��P��D�v��K �'��n :� :�N 3Z��@ 5m+Mh�Q�&@�F��l#L\f�u�pp��)~s	�˰<c�T�`s]&%m����Nž��S���׿{�F�c�}�� ��xB��� ��D��0�)c�0�E�pC0nW�d�:mQ�k#�u�(�L	�3 �&]	0n#ص�d�`�y}B���
|��$dW�5 �O��#
�H�k��%�Ѹ�H��! ��,Gu�a�^(	��Z��{�ߔÖw�ð=:-�F�r-U���&��	�[B��sǸj�8�<w=��ў����cP�jh�{��8 :y����[1,}Ffy`d�z��Fen¸����K5��c~`j�ta���[��_��x�|{��O�_���W��W�S�O*nGӿ>jD�㪽��:�L	�~���8t�a�;��7�x:́��>uOgC�T6�NBOf( :J��<���O�]T���\>�����S�R+�)�˰$��ػh oI�w��� *�╽C�# �����}���E4z_��w���n�][
_��g�������S4^<� �U-�?�X�c�Ւ�UKL�=�R��'���o��3�_ç�ɻ�'�8��X�	��Mhx�8a�7>����7����o��'o��_������~���5��?h���~�_&����~�^�C�W\~��+p�w����0*t�a�Jx���������?�K�^GJO,���8n�d����%����#C+~&F·��+��`�rs�L���+-�5��|�9�%�$mpD�r��3�v~?7M��*�	�\h���n�Y=	>,�������0��:����~,��Yb������VЧ=`k0��Q�	�kl�b��xlu"�:k!`�.�f!z�)b�M$��"�ǎ�����,u;S1��=��#D�1A0��E���_�@�t��:'=�w3�bN�tۃɶ�d�+��03�i3m��I��A �3*<��/<�m�Ƶ��K�f�2�\�sfN���#�&���~",�LaAM�5��abcK'>]��~�,���L���d+�N5�զp�Y�ĕp�Z�>d�e��̋��⛏��k�q�b��sB�`~�F���w^�,Iހ��@��/�� �{�(�[��$p1���`�?v�`>z^S��kJ��$e�o¼�5�L��\�lD�LBl[A.T�%�n'@
d
x
tn,��£LK�J�	�j���b �H��x+�2��/ �A��ڕ��v�l��v�(í(� h ���U���)P��hM(<+�UtB���)�׿˯���OI�t��+��7�V��l�֗o�gc R��"�b92i7'�F�a��!��HH ���' )Ig�G�K%��/&��gO��I�-!��ƶA�3��s�����*�@��&AE 4Y2��.U�O��3Y2��A��,�cL�)�)�<		M9�ux�d�)a�{�2�~br�U�U�
|ʴd� �a$��÷( J) J0�:u£8���ʱ�#(�$�y7 U<�}XՒ�cU�%�
���ي-+�#O� h6�>��9M�����*ó�C�%Yū+�
OV�&+Ӭ�_��6sxd@ߔ���ĥ�9I?V���%öH����f�z��w�Q�)� z7 ����>Y��5
�@�w�#~W:��!���>Q���t�%���
|����!�3��)©��q�qH�]. Z�E.�ߩк���p3v���R%�	�"�К�k	�5��P�r�[��z�8]�,>h�|�$�v��P	ŕ��2��24����:��x��=����3�(��' M�K�w��RJ��Q��"Њ+�8~�"
��j�5�ѽz�:��d+GK8Lv��TW����w?����������	����BXB1rjQּ�=(�ه��f���/,>�|���S���T�����!H�.Bum:�:p��<�Ѓ���u��՗�/�J6�*�A����U�'�~�gS=ď_�׮��g����qt�^���AW'�كΝ�/��/?�?��-�+�~��X�CBw%$w P����/���Bi�B���z�,^0	�Q�����Y���`���b������x
��;�}��/����v�9*$@�'h�h`�vɽ�����,<S�{)���^�ERC���Z�kKG"���ږ�xI����6.llJC8 ��5qH�����(�S�ە��^~d��^�@�oI0�P�̳��q�( �������� :z�hN���9�M�A�F:4:��t�?]F�Ma��6���9�Bcq�:�#0m��j6j�Pͭ3��6��\��^ë߼��?���XD��y�7ꂡ%!��� ��+���PP�j��a|[4[#��g��Q�&p�T��6F��bA �P��R_h{A�.T�vJ�[�}I�X����`Ώ��>�PL���Ʋ^�@a4��0�=� �{	�#9�!y�j�;��Y��� ��Q��K�A�L�g��:+6�Tz l��6�������a�tw����k��c�A����[}<��%c}S.�;���S��Zl���J�wW§�;���Z
���k�1� ��s��|=��b�6<v�I|����K�i	�����D�R��WK�;�����[���N�����/�������~���ą��7�� �z+��3K�:�jx":���Ei<uN��� ��|��!w�O�0�M��C(e^��uwJ�R�$u0��x:Ҥ��R@O���>���7�;u�� *�ܹ��������
l��uK<�m��T$��H��@	��-	�����{ԗ��|~7�m@�K��?>Ż��o?�10�V�o��5�'ڻ�`��h��^Ec/�L��� ��(!��A�.��8OX�D��>\��s�S��w?�z��|���_p�w��[}��}%a��|�����|�^��:�����{^����<������֙[�M�����@��W~�߾�����
E/�F�jO[�����)�0� :2z>���w:����at��,2��f�.@n�|�m������
�s��}t
�Q���o�#�.����X9��Xc>�s�8� ƶ�`���fp�c;gC���νp4����FK(�T��A�κ�l����Rd�P�h�Lc��0T<���t:E���w�D�4}q��z�ꪋM�zX笇5���.X�j����eM���I�`g�K��pu3���㏠POl۾!���%Ly�c���X�f֮Z�kWb��Ř6���e�-a뤒�$XM2���,(Wk8�pT ���
�&��A�f�Ʉ����vɫᘽ�9�����<q������c8|���� � �Wb^���ߊ���X���;�p���x��3���A��������������������ՑX���c6`N�*� �Z�M����׮JB�!�;5�n&`n |�'<�=�R���m�GI�����Ty>�o����T 4���uey��uQJ�L��U��2/�)a����IX��X8/u�U�w�*��W ���M�t/�Ɔ��
tJ) �6�]��T�g� �Q�x@=��$<����l{��L��8� ��o���I�$J)�O)�	Y2&� N���?Q�\�eAS�%[��P��<���[)C�.i_>4R�xDY
$e�$lWIT�}H���(R��JX+��mC��J�F	-�	x��;*a����	l�=�����IN��S��n'�+P%��� T�jȔP[9w���dIB�sUO�)G�����҄��J������j@�:%L��f��-P ��B���9B��uO�xDU�Ty����@S)�p|*}Gy��O0V2!+���4����t��@w���z @	���ci�p,;��:�@g��,�MOw�@(�2�7U�&��#�PZ�U����5JF�����x��+�pe�"�P�
^4Y��?��T�BЬ���YO��0���)I�@:�1@�@�=��_��=O�GŉjԜ�C�Iɂ�� *������O J`I�AQ�J��#g_\6��^�{0�dl&[a�TG8N�\',X�W
_��;�w���������\����iB����X���K�F|^�2�QN.�Od6<C�����$�� 6�QqHHLBaA:Z[q��Q<v�A���Sx��5|������o�?Һ�y)�Z����~�/���"��w?��_��K@�O���k�c�|��W�����x���p�ū����������p'* �C��*�X�����;޺�:a3'��#W@Nf��ع:�c	aT<�'���?|����
>r{��b�>܋�˻���T	�N�_�
�G ���x�%�:����+�Z�r���&@���$ �%1l0B�X�U����Y?�f�G �,I�IHoNG_���4d�f!�+�=��KG���*T<������m�x@����������#d�t�t�u�KCĐ��l#/2��j;�mv���4�
[��l�7���V�ul��ܧcCE:����w�ǋ�^�hdC�ab�'��� ��PP��PEPM�NGt:#1�=ZmQ�m����>��~2��Yև��皰�+��A3c!4��9wo2>d�j?E �:�s:�ラГqCi(����v§��@G7�a�x�j�oR���1=��3��y� �/Aѥc�q�$*;���B��b���p��gp���q�Ƌ8��K(�w���!ƻh�go���x��U<G3��>��_�7~�
o��#��Ox����O�F}Dh{��7�������}����e��>����m(:����f�|�������#�/_�@@yO�%���_g�+�~�����?�z�u���,��傻*�� �#���k<x������ޓ��l�\O���\t�fC�L&>'F5��x�is,Mz{8Y54aQ��;�� �)"�ԩ��$� 8�y�n�ۥx	}��������T{;o� "K��{V ��A��0����)��P۾�I�Se��]�H�[��;5�����{@��$\C	��rݑ��q$�ҡ���p�o�o��e>���?�镑�����;����=���ͮp�6��m�?�����������#�<N#�sr�`��	�'k�u�}�� ��z�2�|��|�,��1\�q�x �?�K���/�Ե+8q�2�=u-���l/��ۋ��w#t��(�N�vXW�cFu(���o�$�������`�Ʈ�e�he����
|ޓ���`p�hE/�9��|�,�Y�e�f/2��U6�D�و������\b�z��C��ƚIZX9I+]d=,t��7�,̧�O��i����]��еӄ�S�M6������� �k���(L1��L-̷��r�1Xe5��&`���rߞ<�����~[_7]x�hc���O� O]xp�f���E<��OC,w��bG]§f��b��8�����\��h�+���!:6a���شe�l\�Mk�f�b��֯Y��+�FWaղ�p�dks@'������.ְu�Rd�F؞b����N����5,\-aG 5�l	�)a�n*&*]�6�)w&e��k�"�����L3����tm�,d�aM�;dnƬ�M������#�,���ƕ��p���(jI'�·��ɘ����1v	�r%yњB?�6@�:'tE�YZ���TB]���,����*�)�)�)R(�p���TP|��,C��ke9�p�C*`*�U���M� �m����a���TBl)�M�2��y�Cs=�.
p�)�Zn/��7�*���@�^P�P�w���P��>�B��8E:����&&��̰"IF��L�z&�U���g�x�8-�Yp��*����S@G<o9өF�!񾩇��i	�og�%q�(Wϸ=����T��X�y'$�n�*�T�I�&��˲y�4B]�%�l���T������Q<���p�r��I�T{@E��x�N��
|Fsۨ>��n.#�JX�Pu���a��JWe�n��S��=���5+*��7T�C��~�
|
$Sj �鸽��u�̷̑�6r�����y�J����m ��cd�}幉d(	�/�x@������QOV�a[Qy� �[���B��>�m��ܙ����w2	]�
x��}&|�>Szӑ��zY֓�^�ޣ��8d�����=��1���%�o�c2Kv>P��5�� �&����B��T
��"��R5��T���m�N<$c�����ؠ�����#x������^*E���� �LTRA�@K�e��C�Hߝ�šK0�a4�5`�2�.�p���s�`��eh�ۍO��vv�#<�]^�c�W�̪>D�6`sD6�E�#��E�'��xI=H,���\l͆oB)���T��*��'�'$�i��/AIi���QWS��:��{{[p��)�w�:���c|���+i�������駟�ǟ~B��^a�j9��W�����J��	?}��EH���/���7y�7���o�Ox�/���?��?�>cܑ�����T<�_�)~��ط��Y���`�f����O�o�"�������u����\v_�D��|�*P|FRw<d�=W��I�r	�ҏW�	�Jn&�W{F՞P@������x$6�#�F��רT�Uӻ4X�WE+Ʌ$�P:�S��LUI�!QZ#?n%����Q��
���0W��9�t���@G@�q�p�����/z��a0��˭`��.4��������X�)��/�ٸm��;�p���� h��q��x����荧�ؒ���0���J������
�Vs0�7�+}B�[	��J��N;ᓠi�=~��z���0ٗݦL��%��q���q��w���}=��l��wE)}?��B���%Ö�ْ���4h���poQ�n@��a\S0k��i��_?ĵ_�����R��(�����W���������������?R���*_8����0��Q�fx���9e�
	FU���pUU�o���)���7����? oY�S�a��l,�3��)�'*�v�����R��������������<�*�/%�``���7pE�+K��g��T���o���%�+�}YS�r���/�y]���A(���4,fC0����\X�ɅT��ީ����cI�N�E�	� `�� ���N�!T���T��� �
p��#$JB���$�G�g @�H�!	��&B����n��O,�Vo��>)�]��[�@��[o�n�/C>�(���=s��5&��P2Nk6������]�|�A�-5��������XޗQ�F���PK�wi�D��Z��W+in�����4��I���8���M] �	��J���!
��°zg$�UauE |�џ�о,l����GS2|;���&r}��( ��a���a_��� X�* ���w���'���/���7P��
�R��)�߲�u��
CSV`�(q)�$.è�0�^
���0]� �eV���3�`�:'�OE�&7DntE�rl�����^� ��e,e���#0�r,f�f��M3�t78;�u�DX�~�R�r�-5�o6zF�`�?�Z�a�1zc1i�.�Z�a��x,�8��b	�_a�Ii`������-©&��h`��6�iT��������l����\d�s����4k-�Z���\v'�Ŏ�9��� $�������6����+xVb�S�S�Ĭ]�[6�V��ّPin�I6p�b'�q�����^r]Ls��;X�����u�`���p�1'N���4�r��#�j��11z���:}3���7ƃWO�~w9��>���aF�8�/Ü�U,Fۇ�<����CQk-���ď]�iI�0;k��p_��I�0q�F�%��%�.Ǽ�eX���o"�h �q;!o+�N��V_��ɼ;�ӣ2�E/�s;|
<J���x;@U���(��������:ӕ\YOBnUC���S��H��S�����>)�Iը$a��I=K\'�)޵��[�U	� ��ܭ���|��� ��g�1�M�	?���y�
�
��b��[�@��U��R-v\�U�
t*"�(��x�8,EE��'�@I�C M��&^Bt9�A^�=U���e�Ѹ��R��<��D@M�'^RY�2#��|[�'�)!��~�wz>��;B��)B�O�7TJ�2
�	�)�~���2'�#ɑ����S<�"�z�'T�����z�N	��~��
��<�3�"�l#�$&��od�PIV�LV�e*�:��H��DQr�x<�N��3��)`*�R*0? ������!ZR$���)�-a�"���4��q��f�oD����V����D��q����ѻ�'����v"�6�$#J�#��dB��ihrO2m�X䱮aO9z� �K�h��KIB���N�<��Ӎh|�	;)���Dkh�Ć���$I����$xʐ+��S�W��Jn�����|j���k���<��s���!�VIB$}@�Η"�l�O	|J�.�@e�B�@(�@��|�@D� ��&󊷌�Rt����£%ؚ���l0�j4tl4�A6Ǥ�p��YK� )7����6�E"0!����mĶ�B�d�|;�������Eq�)�^���G���]Ҏ��E����
l�.�{d1���as8_��
��u��m7��������X���{�&ą ')���h�Y�}�8}����!���ￋ�Ee��A-a������7%+���O��S���W�rR��L	��|�)>��=�}�5�������w�ѻ7�³�⾋'p����/	���{��;o^�ī/����������#~��s6<'�{�	�v��|Jϕ��th�G�8���	��g�Pt�\�*���r_�TBq��w&"�9��IH�4�B�×���#ea��B4�ĺD��)a��T�$#�R	�q|��KÕ܈�XD���l:t���
�>j8�D�*��eX���1�Y?�Y?T� j�	]W#�O7��3�-���Z�lq���L�a���3��HR6�h�:ƭè5N�ܙ��o>����|��*2zJa�F�[�W��:h��cB�/���b\�����M��3 ������>� �mɊ+}6�ba��bo��/�c?��$/y�:�٫X�k�S���d�ʂ��,��fʏ�́ذ񓾠���#�;B1�3�ۃ1�]5D���w_%���e������OD�Q?���?��������w|¨?���կ��?~�)���;��^��=T<ysZ�ǆzb�����'/⣟>�o��W_y׮=����7>����+,_Ǉ_��/����^�|x�]|��Wx��p�בy�S�|�����7�l��.w���to��S�x������o��߿����'��7�;)}��zu�*��H�ʢ_	ìS�m��;�DG�.IƸB��Z|�޸�"_ڇ�=l�����{��r$�ǳa~2F�秲`x4���L��Ä�#�|$#&*�Q��$���%D�4��C�L�2?�_��U�}�	��)��:wzպ�7���n ��>�M��<��*P������-)�l��6	p�����="��e<�;$a���r�wh������;��r-o��k=j��OR�
L�#aX��v[���10���;�#��c������B���C 5�!�6`h�:�^��a�N(폂��F�7�����E�0��b|�h�.�q�
�n�S�V8�n�C���xa�a���\����Z �
/�Ux`b�7&����aK�5M^���~8��Y|�ˇx���x���Pz�S�`v�L��14i9)Z�{���й<a�a�>cg�C�6L'kb�\c�Xb	��N�<�k&�c��N��R;,$p.%����E���Eg�Qp&8:YN������ho������N�!p��.���@wt'��6��v�ڊ7t��&���i&�0k�x�&���1�p�s'�Q4�Z`<K�'`��.�� K��� �mu0�Z�<���X�r���6,'�X`�{�|l#tnټk�,%��d�l�X9� ��7�$�
x.ƺ�K��|�\,�?���`��=!�����NWع����N3&�~�t�#�/����c�ҙPk��x@M}gC/x6t�f�$rL=]�,i:.���w���܏��������]��g"}&@'�-�{�v�v���N�����+�cA�2l(����@��v��6W�\`g.��}�!|�[��a+�d��S�"rgm�J��ņ|O¦*ѐ��)*�)^�;�x8�v+�!���Z�UK�S�|
�&u��O��%�FB%W���vY�ݞ�H���Wɂ�} ��[M�l�T�|� �\��hU=��}@LU �@�Z�#�v+����ro�-u�VBh̾@�*}@:B��~��{	7	��Cn%� �ԉG��L��W#�'�җ������	|rZ�����GJhoK&�b�b%\.�V����qi'ס�}����v������K��~�ҟ4���]nA��]
�FdT�銤��xB�s'Ys�N�3�+IQXO�i��d�U��T�U{B �~����MeZ�+�L�M	E>J@���u�����$b�6
l*�)�T}B�u��[�Q����E(�>�i�
	��W�N�5ZΟ����	�
��Z T ] 4~7�U������8��M'��q�0<G۪�Ϫx[��5���M0HB�|������>U��X�����@DC<bZR�L�q]�J?Pu(nro��)=����^.�L@R{���nw�jК�vb���)C�\�G��U.%Yp�.In����������vT�oB͹fԞم�M�8T���V tϓPu�NIB��4!� �I�n��*�q!�����PG�nx���M��t� -[XO����̏��E3�z�&t:��G�Nq��.��Ú�4eԠ��\|�#���Bx�.��t^D�!���y�؞P�M�EX����[���u�@jm��]AC'�v����Q���@TH(���P]T�oOzlCD�2��P]���x������/i�
l�A��$Ң�i�*�$(�����7x���8s��w�!&��7.��-�8���2<��#����/s}�
����'�~��<��Y���nᇧ�\v�݁����>��y���.��O���[���"?���и���eK�LFJk"o�Ҹ�~K��_� �@�Y���X����g^w�-I_PY\�ƣX 4�����k� �Q*�����0��0B�p>�a�ǰ�������z��a�C���s��/�Qٺ�a��L^��Q˱(n�emǦ"?x	�V�!fƮu�7������_�˟\��o=����D��Q�T@����?B5(͆ h7C��_��F��#��[}J��W�� J 5�ɪ=&l��ƣ_W2a��۷8w�*VW%cb��{�`M����w���|�}iJ?P���J��]����m��gW ƴ�¨#vDH<w�i����v�i���#x�ͫx���p�����k�W���O�7�#���������W��o=�>��3�<�(~K�j��[a����\��	����x���p�sx����҃���}x��\��(��~/�t���W_z�|�~��;|��7�����W��F��]�����{Rt�Yg�Q{_'jO�{w�{����c'p��Gq�W���_-ePI�%���G�4�����{�������O���_�$�,'t+}L�éd�h �?�����u<�c��z�����4�ֳ�s �aq"&�O��ީL�s���Ɖ�hL��C�z8E�R T�P2D�}:���,Q'&��	x��y�����w��D�k�m��+l�M�o���B%�V���k�xKy9/�{$��8"H�5K�|04[ ���q��ݣi�ޟ��|��^[B�;��~��{�0�3��X���To F��ch�Fwbt#˚�W�Z�0����@��=uh��m�lXNi����XL����(��u�q\�8vF¦3�a0o�Q] ��}a��k+�p�ɯ��/�ї�ǎ}XH`�U��4�'�lǄ�����bP�"�X���sa��!`���f�A�j;�3�OĒ�i�<V9`�R[l�mF���\��Xl����L¡��H8����HX����x���`gk}��,Ez�LԂ�DXۚ���f�z0�[#�����DN�ƙۻ���+at��xL%�N#xNS`��`%���)���	���ڰ���DB��,1y�,����`�֕p�DP[�+������1�Z�p:as֬\����s�\�Y�+�JܙX8o��r���Θ6u��8(^�IS��0� J9N����5̝���ES1�B�[36�a0�J�~s`��`5O�
��'<v�ׁg�z�x��a}�̎\��05s=bcN�*$����\;N]ރS�G��JD��Z�m��	k���m��	4E��g`N�:̎X�Y!+0;d9B�*IOr�"�!��d�U��JOu�!�л(%ɄT	�RBo>D�Ą\GBqE�2ơx>��Ӕ�C���Ͽ�����V�rJ�[¨���i��J�P%!�}*�I�-T��)c�B�IV\�����W T�lT �|���$DA�!G�d��3���H�	7�m�dFM�+����� �*3�x�ĆVyB%W2�* *!��9��S{��d�l����f݁,��Y�ʐN -��@;�� [Am�~�H����J	_oAT��V���>�z�G�o�#��LBUïdxDU���}?%W<�
|�!�OR�U�]*�'OU""��74^~�����$P+^�P�Ϫ�� �Z
d
\JP�2��E T��T��Ǌ�5��=#CNV ���p*C���0-{x��x��x8/'��@�x��T���*p� ��{ә��]ш�JT T	K��C{T ٕ�ާ�+�h:ۦ hq2;w �1�������U��F��u��+o�Ӕ�
��@��ܑH;;]	�U<��4�PIB�d�}���0,��I"����� ���� ���͗���@'�.���@Z}�	U�Q}�QIB$ *!��-;IP��P^P�PE���{����*<S��'ڐܙ�A�a0]_�8��NN30w�l�_���Q��؈��n���Fe�a������|�W#�a/���#��J�G��Q�%A��L+EX�N�7�?��r��/�S+Q��>�]xqU��H.BTa
{Q�ԃ�xx�"-9�����{ ć��������mkCnz*j�v��=x�+�q�5��ӷ�c��?����Іjq�O�F�����p�0[F"B�=�+1o�LekCm̝9A~�(/فW_��?Q�������_����cߥ]h�sSs�%���'� �	���@�$�)���	���+��T 4�5NP	�����$ *��k��"E"�,�lCJ�S���,dv� �#9�yHk�D8(�� �)!�	�4�9*!��t���\~EP��� t�(��u��A���s�0q�&����z�V��LL]�q��,i6�y����O}6U��)nƭs�;�oߋ�w^�K�F {
�텰_	c�QU 4+}�"_h��A��_�� I@��	,���a|=T��Q+���Z��aV���x=@��a��M[�J�A#��w^��?�7��'���������+?<6|����*��=��aW�H��<�-C�0�9 �Z��舀	�ZP���8N|����Գ�����s�M'��8Q����م��(=ۈ��,�P~v��4��t�/�"�\#V��o
��N�E��;>~��1^}�y\y���v��@R��8Y�ܳH>]��}lT�������?�'�|�7��|�>.�"��a&�ֶ-n]1�ם��lĢ�T#��](�ЌR~�v^h��G������īWp�g���ޗ��ï��;�&>�����-|��kx�������ׯ���.���~o��>�����R���%����^��<��#8x�8j/tШ�Fܑ
�X��uw쏤��X
�OfB�d�)��:��#��7T� :�̨���?�/ ݟ� :�@4b_<�K���*)�$W�OY�uR*0%����@�X�C�zC�]=��t���x��*`�]��Q��ީ�_�^�����@��!��H.E"�I�wy0��dD2/P*ゎ���hn3�ی�6#X��~�q���]A�JHm���ptW$�w�c$A^���'#v�r���v~�����1!�N��{���>f}�p�;�׊ǰ%��K�[��K�4>#n{����u�aMY���	�f|',����M�6loNţ���/���s��tj��ay�F̒���ް��Q��N]���Јy�Cga���F/�Y��Zd��3t�7]�s�1k�	/0Ú�V�L ݼ�k��b��;�a��x4���^��F`�����Fc"a��TF��)>Y�gL�h�Ԅ��V�^�U���DLd�)�5�rs]ؘ$'j��L��MGj��6�,u�lc�I��]XZh��bL,���oE�ф�#�1�+=�!(�ۃ6b����o�6��شvV-����1o�$,����<�LS�t��)X�d6�.���9�\1}�#&������S	��Ӏ&>�j�fkB��g�Z>�-T��΋�b�<���c�Y0_ ��0����^np��c�xJ�`��y��E{�3`v�FL!�ZG���Bo�}�8��a�Ѓ����|��%�C��Ya�{g�c�4-�m��,0�k>fF�ƌ���3��`n�R�N܌@��Y��F0t/!p�ϧd�Ug� U{Bo�vJ�R�t
8�T���˼ ���
�
�*��&+�N�*뫓��T���x9Ua��F	í�U��W�s�+�)!å~�ˠ[ *��/�x>wF*��˹�PI4$��J<tw �T�?����
�}�P� (A������-q�T��R	&�T T��V�`���d$)�$�
P���-�'t*0J) J�R@�eaL���l
ϱU�m˱��N�M�DDф��>�*	��=�(E�MIfݣ�(��,/v�� A�K�aS�S-�E�S�%W��*�S��=�[���hXo�\�~��>��w���~��/ z'|�M����4�F��DD��	ܷzh������WBr�U�w��G�Q��kI��H�=S�"����%�@�L�c���� 4�/	�i���m,�/�A�t^���8+��'�b��v��Ӧ�*WBp�Tu@�hTs"�Zݞ�xA%7Q��@�h*!8�=emyP�a���/� h��:e���� ���)�p�4������;�����S�� T����l��@6��)  U���@b$�=M�4��T9�
�`Ǐ���0b�e:�γ0u���ÿ�c#��<���|�7>��]���潈/م̺=H��F��~��?O�CN�!��v �����H�oGLy=b�jᗙ�%��p�����Q��4R	�I��(�;���~��`G��콄��:�b�?�x�0��w�KϽ�Kg/"#)�[�����XT���Ⱦ^<���������ן���hU�JoI���r�?�����~�>k���w�=w
��|�#������y`���p�����%��� 9>Μŧ������=��O��K�8�x/���3r�� ZD ��j�w���$��+�P��J&\ɂ+��O *P�Y���e#!�G4���E�
���)�:!��ADM,���ה�h���#�y���:1�	pX�$!5~�_ðP���*��� :� :D ����	���r�,�9*�������?��ca�Z�H݄-����1[k"09i34ֻaMQ:�8�+7��sｌ�_i�E��X��-0���f� |�j��P�(K� �P�4�@gW���"B�NG�Wz�	0h��ec4�s����g�����}�N<u�e)�T��tX�IS�S��Z ���3$ЈGfdK0F�P�+��B1�3\�Ř�kX���|"L]��M���8��$�JU_X���1���}1�d;��7��x�	��y[`I�m�I�'�[h8�%��7c2�aYk*��8>��s|��{x�P�ճ����F�k�;�vl�i�g��[�������x�����7��_�oo���BO���1	�N���^u(^|>c/U��]h|�=O����'��k�����8���W��{�����>�7o>��7�[o?��o?�w�z 7�}7�o�����i���sx彫x��p����^��o���!�p)���Ʋ�d��J�L��<s^��Y�9Lh<����r,!r�Q�G�1�0E�e,t��T�ڛ����0P�ȽKJ���%����@U<��	������n@�@���@u�uu2e|ػJ�T~+ x7PL�,z�`�/t���N	l�1oW��s�w��(�y���U� ��::�#:��H����t$5\�t���!T��v�bd!��'}������!:���p���*���{�	����)
Ľ|G�G`lG��>�h�h�C_�rO",�ba�s2㽷&�����aw<��v�q�ꎆEW&v�Ôۛ�}0o	�5�V4�mr�c����~��x�g�������N,MZפe�)����1!}F'.������L� O��	��Y��6c�X`���:���TmL������l�D��o���i���c��6�L���h4�G�J4��&:�`�M鎁��8B�Lu5`�G8�׀.�T�xL	���B`�=�v�Q=-�iB� jh��gh4�#��0f)24漕��e_�V:�z�s2�B���>��X�i�4,[�� D��/���[�@u_F ��U��`�4;̝l�yS�0k����S	tΙ��� |N�l�)��p�$�V���N�ä)�p&Ⱥ�v�ԅS1o�<,ް�7.Q4k�|د�
ˍ�a�=��S�1��6���H���0x�v_�B`a�Ƭ�Ԕ՘�o�|�Ѷ�0���zo�*Q�Y���p���؏�=n�>o"F/���R{�/��ɾK1-l�>��/�T����H�ų0�{
h�&a+��u��
xJ�[)F� z��S���S�S�U��:��TyHe����v\��v��4�V��HBtUI�T��*$������T�sنm/#��'T�S����Ve�h�N�>\�J"Ʉ��m��ުu7 ��6] 4�@ᓶљb@U�O��4�;* ��%�SU(���;�GR�ӆ�tN�'P�%�PUU�	���������6��B�x;���#���U{=�/�$#����OT�#���D���_�rLII`�d)^Nh�$�)O�P�* K`�e��C�j��L|ʴ �:�O�n	�%��o�]j UK���Oe�P�����k4��yI��)`)�j@U���W�z}��uU�K_N�K��P%�0��$i����+��)�O �Г����LT���vRtP	I��Mh�Ch[�����rN6�xw���+�?C�b�[F[:�u��	����H�kP8�@S	�i]�J��]٪,���H�2讇T�����3�o T=6��{~j.P!���[P���>���x}O�C�J��+�W�� T�>\��w��r?ǲ����Rj��2h4��Z	M'6@�z0'�̶���Ip���k���o|�)|�j��+�ǫ�ĮC���ch9��O?���s(�>����#7?ÅW�D���Q�gR�k�������GM�!�t�#��aUέĦ�,,���Ï���?�������������Ĥ�q���~���"35��mF���ҊDd'F� -;+q�@�t
/>q�__}���>}���s��S�Ȱ��?dZ����ǅK���ڊ��
�壺|J
s��Mشn5!���ʀ�{�����p�B/�څSv�$��b5�.���\	
N�9&I��EU��#�[����TYp�@��E5E�	G +�"��q�)�"�Y� ��?l����|_x��,T�o)�� �~K�6g{"�<�1��1�0b�0%�n}@��C	��j��p��	̗8�z��N�$�p���y��� ��"?xW�!����LN���S�:?m�����=��n<�+�<���b8Ƭ��d����h<�$�N��K?�ے	�j��ns��� ��͎(���+jE 5����8��u���p���q���Q���`8w�(�@-���bo��k(ó������F�i�ؖ�k��NS ��kTm�8��c���������㇕�R/$l�Vn�c�68Tz`R�7,j<1�����0���V�v���om�&!W�Ʊ�n��vL�v,�����O��?��W������bLJ� [B��mT��M>0l�i]�2����\~�1|��w�?���C�C�1�4�-�ʸ��4ʍ�"a�
���h��Ec�C�� �\Z.7��J�<ډ��;p�^�� z�8�|�4�|�$�{���� �����!!��+x�z��K8��^t�mD��r�Q�GkPp�>}��ԓ�%|槳aq�I����t	�.T�������={,c��`����~��$�m:FbICet$�n :r_��VR��rB��C��ч��R��Nϟ�v�T�����x<o�@��pJ����M>��	 %8��-�T��W�S����s3R��R��#�ưO����u�%}�)>wJR��`i��UW��r��<ν|'���1�9 �	��Yi'�F`d{$!6C���z:	�|w&��5 ���ab_�	�VOʲ��2싔������5��xg#1�P��8�_��/��ϼr�9��CX��� ��E`V�ƹk���RVb�sx�|	��A>����#|'C?`���3�c'����hX;����̞���2��L3��e�%.&�i�����h���F�\w�����D�ШGH��	��5���	�㠫7�J�$��N��U������D=EZ�ژ`�A����8L����=�4�b��P�4��+-�F0�i�%�0_��Z7غτ�?�/n3�Gn�Ƹm�K�W�;ܽVb�֥غ~�@M��<W̛b�x7�2�tu�����N�6 e��l&Y(ð�9[�����s�鄩�`�ҙ
�.\�K6/�r��X�3�-���BX·A�\X���}�
�M_����r���� N�;���N��%�K��]4��!�TB�H�PrU��rP�3�c�C{�!F���`<�s�"h�z�p���bL	Y7��p�Y�)��1�o�.��,/�wd �9�;��&o��y@%W�|��aX*&�LJ�H�멪�T��!�R��E��x\��)ö(�I�TK�S=���7t�N�4eE��	U'"���� �^�O��R�SBq�?�� T�z�]�ޗ�����J[�����3鴑dl|�	�(�)���U{HeI�J_H�����_}$%D�� �x0y\J�T�����J�PIT�;�X*}:�8<�l+Ʌ�yK	���y	�Uy<U!�j8U��r��=�,���S�Jڄ���z��n�K(+�S����oy@U������OQ�S�@� (�/I�� d�aR��y<�xB�`)�۝��=ҿV�9����P����{��PUvb5�J����n *Yp�^�JS�����Z)׀`Ex ��J`l$�I�����0,)-�4�:�;�F�J��>��)���&��@����J ��LS �}w=U*�I�l�v��*�J�Ϛ�Pu*je�g�Qt���}��?�e4��e,P�́�[%W40/}B@k/��z >kN4��[q��)���+�C �q�ż�;h4��:͋��Be@�	�i|�R	�)�d§J�NJ�9J:��DJʤ����òM�U`4Y����Eh�ܤ�^	�.�v� cW=�̷��[L^�����dMWvAm�	���F��Gp��{���5t��<�/<��O���Z�4z/<��B��(mۅ��*�d���!�{�y��ݍ����;��G`��P�d�BQ�ĥ�wH6y��+0	k7a��-X��i�E��lBrb�=�7^{=���V#,�u���U���RjN;�s'��'q����_�V�2B�������ҵWp��9�8}}{�����--(.݁��L465���6�����O�����ԍ��c����`+��k@��2��-E���B��G�d�%X�]��1 ���?"�3+p9-u�G�����v%"tg8�*�E^ؚ�$�$�z�K6<6;��E�ܘ�hS��	�ۊ�����|6j��e�=�!�AlP�ʢn��Q�	�λ&!�T��(� ;����4vfY�~��6P2.��4������KR�cM�6l.��g��9�QpK\mn�2'm�#＄W�x��Rڋ��&i`�FK����Ԁ'T��j�:��M��R 4D���R�$Ң1��Ű-�Q0���*\��M|��q��/q����S�W^;7B�U2l���0�1?�"0BBn	u�v>�1�5�� ��r��5��q�g�	���|�w����0�p���a��4��$�yw2,z�}a0��mD�]���ݑ��V���a}~T'�x`Q[*������|��Gx���]�������q�/tZ}�Gcݐ�`�B0/܊�襱���7q��x�7P}�޴9&ݱ0����ǐ�O,Z����94з�G����}��t6;.J�I3�����J;����'����~�?��O����6TܷY'��F$`w:���cSk,V��Æl�8�ѵ#<ZH�١LɆ��\˃����{�q<�B%+�(�8��9�`�R������x6� �@&�S@T T	��n,�5\�����Kب�S'a���	�wH�Q����8����T���c0�pA��%a������{CCT`x��T`�N�8]6N�(���."�ɲ[���=����)�d_�rY��]�r�HMӻ�.�u)�!R�*�)*	��*��(^��ɔ����Q������p))�*u�����9��:D�%�6�:1�=������q���P����cZB`�G��Ob)��#a�AȌ�}o"(>�V���d�5�3[������0n�Kk4�Ӹ^_�#/_�ǿ}��׮���(۳˓�c�ƺ`#��7�8tr�`|�
O\�{�faP�T
p� �I��ۉ:��s��e2�Y@�UF�����cl�\1����0�R�5ao4VD3�0��9t"A�DgL���Xg,�t�uz�c���'��s[=C������c��q�ӱV:�Kh8�mt`�l��n0q��Yv0�7~�dc�ͷ���n��:���a�m��S3a�7��1#����	AAp�Z�U��a��<�Y3K8b�+B�fN���I�8�L���)�ma�h�I�pp6S�-�a����Na�zK��.�p �:�r$��bβ�X�nVlY�u��51�0/j�%l�|�?����)˃���b�*���1�Ћ�5Hߙ���h%Bg~�6�H݈�+�(b5�2qߓp����O�']��j�UN��Ö�`�2{�_b�5�Рep�]�p�)��0/t�p_�?f��M�^�P��%>X�v}C�/6J7���&�K�\��8���~ �1T��6�¿���6տ� �s��&rޗ0*���Z���xG)���z�M׽�[
��Nݾ��@(�G��� JKEҽd���wM<��IyU�mR$���H���*UH�_�$�~ش���๾��h����Z�ϝ<6��h~����>;E`9��dڻ��a�)h!&�D)r��R��rJ'a,yOס-5 Y2ޥdwU��x�
��F8F @��+�$D"IJ$I�$�V�� �ߓ�h �H`3V��J�9B��d'�1<���l�Kr���,��Jh�2�
�&��`-��lU}B:��j�u������O(�ߝ����z�"S����#�۟MP�9P
�RI���H�f*IQ�C�$�wH6��C���jd[J��*}h�����@B��"�	���g���*(ФM,��uټ��<�WJ���$Ҿ��I�)�cB:�)9[�֧{��D'��z;.�*}M�	���~��H�ui�҅���(#���!Y �)!5q*��"ј�Ȗ$D�%!���M���P�J%rZɀ+c�JXnw24� ����T�d��`;��\��#|6>Q� �ZC �z�`I -��/В3���
�+E6�,^��#�(=J��@Oq����J2�s�
|�>�/�L[	�m�=т�3�8J }�����~��'JPvf
����G�	��I^t�i�T*�(���0�l������q�r	0Y���č4�:��C��"�I H�҇���[�y�-�����f�y�!&7�� /}�y�}T��FJyJZO���4�=���O���ET�=�Ҟ(n�AyG7��Z�s�0z�i�}�A�w�<p�U$��bud4<�rQR��l�~�)t~%�ǑQ�1���ͪA\f��'`��͘<s6nDIY#�sʐ�����"",�V,������(�.�bJR�"�QQV���&��4���N\�����>��m���o��@h�o��/��
|�1n�|�^{z�N�FϾ�h��F���hjkAT|2r2�����c�C]��ƴx��G��ٔ?(�.A��"§x@ ��]�S�(��)J�T<��L�V���"u��L����!�^�ͅؘG�+��66T�v�c^��ƃV�VgnŚ�mX���r�q��T$�R�Z�e\.���pXϱQ�Ȼ�0J�r���*���q�0j�,���u�t8lr���4���Ĵ���C�\���36a]�缝����(l�A79q4�N�@t?v�|r���}�9$��>j����d�4J�rOL �*a����m�.,-���J��^k�UI�%ى�$?i%������I�7����Чo�3��w��_
~u���4Bm$��H��&¨7#h����MP�踶h�e�|���a�cX�a[_��xo��.���<��H�/�d�׆��˂c{
�Ra�K��d�ݽ��R������N�Xh��C�;�E[��9n>�׾{7������؞"X�6���5��VW �w�S�4̵�=�J#�啳x����O⡷GR_	��y�zg��2�M�����<f$t	�ڄ
-������ צ@L#�/"���O�&��6>�^l��`x����Fڝ����&�/m�Ţ�X,��?�'�yo\		.<���X��fv(�46�	�F�| �a�o���L�H���te�ɱ�Q�����S����p��lʲ;��O���T �����}]�+�@���w��	��jݾ�H��T��I ���)L�TO߮{(����p��D2=B�[	u�z�X�m�)���.�Wea5������oa)a�������W��%[���
p*!�N�䵖����]�y	�����)�a�"���v�$W�!m� x`����H��ZN����<��vD�XBڻ��ܗ�d8v%���mg<l:�`���X�4�î#�������L�y�!|����׮��x֧o���Mp(����0$|je��e�<�b�@]1(���8b��=y�a��L��o���2�8MhY����8eO;{=�L2���\,1�L�&ڰ1� �qʐ*j�>M�F��aHR����P����=P�qХt��F��$Ԏ��Ÿ)�Ф��������Va{j��c�պ�21q�t	[:ܠ�����b�V7�D���-�g�?ӣci�:l�ކ%�K0�}*f�u��%�p�c�&��b kg]���*�`3��9�f�auЃ���\��Z�0m-hR:v��sЇ��'���V��Ϲ���t
f-��˧a���X���ay��mj�E��2$�@@s�g{!�=/ĥ���@����b�=F�1� �1d?���ÄP��V��\�U�O��|>'�b��[�a+l1|�=F���ȥ6��urX�%p&��x̓ӶY���U�؛����+`�\�k	dkw�`}�/6��ac�?6��V��2�(�;�њ���x�a8�@�����̋dگ:>�!��`� *���"�o'�n-��|��ď�~�T�S�S��d=�1 �����e�lS<< �k >�����@Xe?,`%$w3�FB�:�:�皢�X��5٦��F(��q��B���J<���c�=©dV������!8�J���e�+Q��O���OۋШd�%|�M�)C�H� ��,K��R4��di�G�~B� �%p��T�o�z	}}��6s &	��x�j �.��FX'!zw.b��BfO*��I �w(F�w�ґ��l��	kJX-�+�`	iJ(1%�/}R�x)��L�RQ��(JBt�m29A�m�x{���i�})�-�	�X/	���; %��V�!%�}���x�>鏩N�rJ\	��� ����S�:�,�����Z�ɴz��%^n��'�U>�%竔�\r���N<�a=�Jа�[�@����4��׾1!��r>�m�G�.^��D^G�^�8�k*�k��% J�����Y����8����h�@[_%U,�����;���N%����֝oC5��L;�O���|7�=s/|�2�>�O�^����w ��Z֑|d�{|o��W��ǻQw_"w��u�+&8���d]LZh���������zBW����-��>�E�H)�AU�u
{|	�^����\E��C�ojArY�z:p������:����E@��/Dxi�:����,N=��Ͼ���Sh��*[��x�>��FtZ9�CӰ�+��z")��U-((�)�Amu�Q�W��GO��e��S3PY^���
��4��a'ʊs������4�W���x�٧��'�����%�:����� ����|�%>��3<���((+�o�?6{nƉ�'�+�}��g��H7z�������(!|*�I���j �V��*y����T��n�#|*�9 �
� �,Oٟ� h@]l��J�t'Tn��|6�%I�>�S�Υi���ҷ�TZ��Y��rE�;VF����YV4Z������7J��P�œ0�}7O���LL��� ]�
��6� tT��4D��u��+3���}x��x�ۏ����#��v��a���;<��
/L��j�@�> j������!iDE�RN �N/�А�����l�)�B����=.�x����V� ���DXB�	�:�������Z�Q�������V\B�D�Y{4,�C��'ϟǓ��w���+�?����H�S��x�M�}���:��0o
�%����M�49��-J��c�E@%�/mM�������zo�6��4�:�ᐽ����~�/�+c�C��L �V�����^=������}_����dX����|h��Ab|W(��p�PZ��	B��z=��N[ � #Ä0n�˶0ش������)ֵ����m�̇2�=1k�9�`bg,۶��2�x<M����0؛�}��ۗ���&D�L��$L8���R0�@F@G�Gh$�r�S��G���v	|JH�=�mJh�x���)��S�����^��;%�e�=�$)���i���p߰�v\��h� �LK��m�GJ	��/4� (�D0	8�"�]���Q�=<�>xI��@�q)ՠ���;���u%ӯ�ߪC��	@o���S<�w�0j����>g
`4���m����� :�Ϥ��8XN�D>3�nvD�����8�>	��N4��hT�t�ƠKW\YNۛ�y{R��)[w���k������w���/��\;V$mƔ�Up+��U�Fg��~�h�-ǈ��5�C�`h��x9a��ms�`'���10~�%FN��(��а]��0!�ZZj��\6fz���+SmX�h���4� 3����XL�����D<�26CC	�m�Q�2-��2G���hb��>4f�Ac�4�;`�"kh,����5.KDng9����{�b�
�����n�.����^ӡ��q�a�����p_;����'�)p��G¶��I�_����[��9V0�e�y6�\h��6J�R���0�m��0�kEYC�9(Ù0�f�����k���k��60�m�k�K��a:,7O��zGhn�}�ɰ
�[����4d�d♗��[=��¦�4q9���%���
#gb��4��[_����~Y�;�cԣ��	���;c�*{_b�	+��SCV) �}�7O����lL@��J�6�bS��bwPi/7���;!T �[����2�3�#a� �׫ T�<��u}*	�ON)��QJ���!ԫ<h R�;J+��2��H@ӛ0)�����D�e�ܖ�)�)���\��e���?(�	��H����@�ig�$��^ T2���@��:���m��Qt�6��Ȧ=��� ҽNl�;�S$�) �s�볔:	����B Mg�ud�	�d*�p�L0(�?��R�
�J� � Q� �|�1��H;^N��#$�#�W�^�x7�R�dN'NS�'� ����$E��W%ԕ���*�+	}�.ڛ�|�L��4=ډ�s��O�#�j��h¬�nta�v�җ�A���c�2�
�@v�.!��3���"��!����G�H/� ��e��2E��L]/P*�z��9�˕:2G$!�j�R�Y��R���e�?܊gZJ-!��{R��<�3E�e���P{l�{���+� ���K��%�������d�_жL�ﮒ�j��W���U �P���V�݅ʓͨ>ق�㻰�L'?u�@�?}e����TBL"/��-,�諸o'��ҬO�̏��ڏ��tC�ΰ����p�7�7�A|��bLY�s�x"*�!i�
�f�������#<��Gh8x��M]��-)CP&�%��D@6�e�N��6�N �s7wv"��Q%�\��ŝ��:���=��ۉܺ�H+mEHr	�o	����LE���x���xq��I$%��駞���-�P<��x��(�߁�x4�7aGn�Â�i|�mF\D(�R�Q_]����>y?�Kӗ4E�O5,����<�����ꩌ!��+�_��7�b��=�x�u|f�d��32q�N�#u���_���*��S�æ"�y8���xAe��C���;v����D6A�P��5ٛ���XK]���v�gsAsa�,���K������Q��=�>90gC�d� %t�Ot��&&�p��y��e
\|f�������bW( ���[$qA�4d���nv�F^6X��}O^ē�\�럽�'�z��E�^�0e�) ZF-'�B5$W����b|�7�U{߂P�E[Bs)-Nk����	O������E�?6���;/�}�KЇ�y�m��Z Ԝ cD��n��� ��I`���0�i�x��{�a�7&]1���}ׅbCo1v_/|�>^��-�{�2�� ����A-"���ۀm-;�|gf6Dþ!��G�<5{��G��f[$�!J��jT��m�8���x��q�w���Gޞ�B��
�T�S���oW 4J��2oj�>�7��_��^��U�t��h\	���	c"�h�O �U��XB�JJ-�K���u�&AR�3�]Q�h�2EC_��ň�Ę`m���1S�e{-§>Aߔ� �i�?���I�ٓ��,���K�ޗ����&c�s�۱/~ <)����B?�U\��� �ZJ�� �?��_R���@(�*��C٧ls;lq��k�����F�r���'3	�	ʱ弤��A��GH!��wvP'����@œ*�a\W�OF���J��@X�J��@<�M���2��jo� ����.����>�%T��R�
��]��"���W<��[�?�h��ؖ h���;��	s>K6���M�u[4��Mp�#�&�M{4&u�c2�t
���}_Lcw����~�0���|��[x��kh9ӊѫ��.y�a��	V9�a���髡��c��cD�L���n�7G���n�ŰM����VXb�<Sh��@�r<�MFC�h���V�	�7���&�05҆���<Y�j�͌4`b8c�>�:�N��k<cL�`��&4�0~�	FϚ��,1b��O#S#�[��s!�e� �>U�ڰ23+]Z�p/Ak��^��1��O���	Z��U��Fs`�Nѫ05v-��W`r�
L_�)�+���~���v�f�tEN��1%p�����B�{q��l�o����`�u,6(7΀��Y����O'�͆�9�^;�˜`���K�`�f*��c�4=���A�51h��JN�`���G�q�ݫ�����ĵ��N�� c��w��[�\�}ո�᫸��#�J���j��x�V�W;`�'�k�6Mg��{!���b���[g��}:�~1�ӱ�d5A2VI̳���=��@K��A ��� hd�&���������d�"����P� ��ӳ,���ou8��oU��>K[e�O�OB�7�5 O�m"񊪼�*��ATRN+��\'�)�-�j��WU�B7��@=	��Q�t����E{+�6t:A4�(���c��=-����G:���>�= ;jCɩJ�*�C;8�@�OPI|sK�Web����*�Z�P�R�q�w��r
d� R��G�S T��J�٬����ۘy��6�~/Bx_�⭋��B=�̞D�f�{��؎�e
R��|rD�}�Ǧ�g+�K��#���.C��*T�!���/�D���hy��D��L.y�C����X���ҧ�@L��������K&Y75��,B��>��W�(H�r���˒lI�ו�ue�O5dJ)���Gu���@���L�^�"���Ku�x�Aa�J}�Je]�^$�˾�*�J�8�Jv]���u�t�dMm��t��ߎ>h��F�uW"����@y�; ��딶g���� z�5�zE��;nB���֞oE�i��V�kF��v�{�0���9�T��PBp+ϗ�� ����&��#��,S�w�����s07h>4�ib��\;�m�+&/���+��=���X����dW� �����ˬALA�^@þ�(�Տ�c�r�<r������Ea�%H�oD����?y�M��ޅ(�o{�D5#��iU}�+iC~�ATv�By�17�Cdf9Vn�Od
�z��7?��У'Ρ��Wz�>v�y%HN������OLCt_��Xd'I¢xD"��!���F\d$��R	����/�?�W������Ͻ�4��s����X��)��S������H�/7��b5�ϖ"�L	�O�t����c|A�?.?�� �v�'S`�*�V]'���S��f��M�<���
�
�Di�������:4+3�47�е9�h4��7b5��9��9/e�mPtk>u=q�G�?|�a1��/ �z@���ZpY=s|�i�T����Ԡ��E# j@��dA�J,I^�UY��$!�ү����(@�Ƭ��bk�L�A��x��p�7���"�� V>�a�
&y��Ɨ�$�����XN�)��$%�aY����S%��15v���NC8��hx�6���k���/�(!�����s�C0��v��st�F�zcT�?l�g��x4iЎ��� BuT��\æP��`ek��<�·x��������?�;?����N��o�G�}�xv����6�<?���	�'h�����;�4�-:	p��͉���x���x������ B��p�C�f�?F�⹉��u%�&��>s7�1��W����=;�A�t�?+�bT/a�`2�0�=c	P�L�ф%�@���N�I��ph�G@�3� *C��8��b��hB�z��O �mƱ�艁�[oo��ٟ�=�N��&�U��4�,5��^�1�1�/Qј�	�w @>���%�r��8.�н]�@��$���G@H<��,@��z�����]$ˆ�z'�K_F�SmO0���d�P��P�`��Tʎ@��K	��/$��y4n�4��\Ix���T�o���,�d�?��稽1�x�	���w;|���^ª:˭x���,��|���$ :�`z{(� �`>g�k����A;����
�e�"�J�R<��ϑ�1��b�N?��������@tF�zo2�v'�i�x@����ܾ=v1�i�R4� ����h�ޝ������!XY�����ݟ��W���z�g۰8f-f%o��/L��������#~���B3~F�����=#='�wk�6S��1� :v�&,���4c�������1�hƛL�x��8��x����8h鏇.�S��a�?�������BGQ�)�{ADi���^��*H���k41&��bz�=�L2�L�w�����c�q�����^\���٧>��k�ǘa��9�Y[:�	��O�z�d�5"�>��)��`���N#��ПE8�c���������=�nkf#�4���y� B
�1.h:,V�@o��W�w��VyAo��#fb�� �nFxWV4�bUS�[�\������h#��o��Z~�H�D��fdh@��Z��6�be�6~ˢ1=m5<��y1&SS�,���Ը%����|c�}�p�Qu�4�k�tiν�j�uaJ�l�
���a4¼	�^0�9N\��X^�i|��p���T���'�t�,�����`6�	!���>�/~x�����X^'�O�9aS��t�d,���!�p����M�������lyv(�v) ����j�����G�dLW��@#�7
�!�3E�M��S`S�2��4K��8�� T���X�T�J�"§���m��SP��)!�*Ϧ@e�R�fHQ�Q%4��)��J;�I�+�Rzӑ<��-�)�t5���Ў8l�( *���s��մ�*�s���o���u�e��O`��ǰ��chy��j�N[�v�@���}�0|�T��:�S K�3�P���	��ǹ>!��T�ٶ�|�R�:@�}���H�z�Ta�����ҟ�@*Ӫd@*���~���M�ܪ�s�`:i�e�W�XF�l�܂��m��
�5O�hG26���=����U�*�@TQV�/Œ������zc޶@�@lm,�y�����\�mI�r�)�6I�#@��� �f�hsʱ����2$��0H�t�S�E����H'��+EAP�GS�R*P8�U�@�:�V���e��#*�Jw6Ur��K��
	��܇���%�U���~$�Q��B��6��x��7u�#k0O�®��P-ð�*Yp�s U�� k��h��4��X�tl�_�ھ"t� mBӵ&4?ւ�! U<�����h���
@[T �N@$"�
��^�A�����v�O��|?��9�����/Go�J�P�ZF -$�
x��P��2�(O�qn�T����Fǝ~�xz ��q�]� }wC8�t��,Wx-��Թ��_���8T�؁ڞ��"����w��u*;��a ��ʐP܈�#а���z�Tӌ��u�h����Z�W5��*�#|v!�g/��ud��BV�n$Vu!���{o�\��N?�>����Wȭ����"���hځ���8{�*�\��=���Uu�ؽ��x��vuc���!)%��Yh��F}o��$oيMk�a]��@�+�c���ؽ{ -�5�k�@kOR���9�R�1+C�y'�¡g��F����~�WೀЩ��y�G �4��I�XB��!)�)�����)��$ :#�<xC *�:���И�X^�Ey+�`�$+J��V 4B���՘��
�	�͙�y���6Bat�F�/���߿P)��� ���<WLG@�|L	�Qh�,�o����I�]NP�P�5�[��3�]���=n.g�aQ�^;���xo~�.�{��t��~�L�$/Ƹ��0���)%���Co���A���F0*c��t���@Mw@;���m+�Zhh@�:�p�ͻx��������>��]��YO�]���(h7��nS4�j��*�A�Z� jLh3#�Yr��~������Ԗ���=�W��	^��u|��ω�?���#��?���+�������O�
6�(�[�jxt% :~_*��Ƴn��F��<L�ˎ�ݙ���u���������"���y����aL�:��,W;6B�,���hx�0���=������g/ u�L�&�Z����P�K�'�{7A�`�C`Ҧ��	����Ps�L�d)�ƽ[���DU%J��J��Q�I�RaJ85h��8�"l�9�������O�'�i��h/�<F�r=¥!�Ӏ�)�'|����j %�h>E�2$��2f�R�J�/��:l`+� I�'|'`�c9�p�����h�
�&�˺;����Qm��$ѹ��2**�G���������s~,��+az"[G�~*`)��m"p�T��RC zL� T$����RϪ΁$e}�'U���6u���S��O��R�6�V���a �� ��X��ZhtQ�P	��i��sH�?[�]��[�?�{���^����w�U��ۙ �#y��2�Fm �ϒl"�ӱ'AP��ɄO�/����ә _����-x�(>��|��÷Ѯ3]���!�ۈiU1�T��L�l�LZe,��� h�L��Z?����a��4WO��`g�X�-xu����DK���j`c;U�O�'\�1���!���`I�=���¨�`��j9��jog:q=syZ�x��O-_k��5#m1b��/!�Bu8Bo�-�b�!�.�G�p�+XS��1��`�wX̛�Q�=a��&�Bw�3F��a�"/L�[��9��({#BJ�U��Ue�"��K_��Ep��Y�Q�JGp�V,/��o��͘��3�C�a1��Σ��!z.c�@gᏱ�߱+	�����y���o�J�J	����*ނ��Ĕ��a�/<��g�r؆L�� O8��N�������{7����œ��c[�6�-r��x1	�����|�$�ݞ�O�����^CD�F����8��M�`譜C�(��<>���@xmX@ ��ߦ�ΏDrO6��4*�<�KB�ڵ
|�@cV�����庖xl�H�ZB⚺M�9s� :�j U��\N`U<���H$���5�	�qӍ�NU�J�M�>s��q=cUê<��2��@&S��Fﱔ6�˲�Wt}g"R%Dt�w�a���FIB�Р�k�Q�t�@����S T��l�%��e8��G��l�ٍ�wv���AT�i˗�>PO(�O�
	�R
x*�W� ���u��BZn�Dۭ>�\jC�c�J)p�}�i{�+[	�M#	p&��V<�J""N�<eZ����74��L%�V�M�L�߁��vc������h>N��Ƕ�MJ\�7������|L`桯h���]�`0q�]��?iY�L�����&���!�bZ��t!�K� mg&J���������PW$����ܗE���d�}d�S�~�$�U	�fA��)Uæ�+)���P 
�J���ڣ�n�!R�^^`S�*Ȕ�(9X�L�����8R��)<׉{����q]	�&<�s�<��-(�Հ�Ρ>��C Z�-��$PI��g4} ��"�S�>�����wC�]��Ш�$޿f%��f+�C�J]��W� -;]���X�C����4�;��ϵ�t� {^�-�������+��}h:Յ��;�S�?��w���X%j�T��J���kF 9͓( �R�3��%�I��8���e��(���*Uu�7mDe؜S����e�*�t9��ՠ��}JV� ��(����[�+\f��m._�g�?h>RJq���y�6�����/��g���[���n'�z�^�5�ؐ[��2�8���1���A�e'���Ѳ��vl�i������GjK/���׹���q��7��7����D��h;|u�G�[߅ܚvdV�S���"n<uO��S'0�/v���ڭǕ�=?��SԷ6�h{At3�n�Cnz&vT{�P\X��m۰-!�i)ذi=bbcPTV��;�е�8�e�"�p3"R��Ŷ�$^��8��q�ً�m�_���b�)_Z��ʑ{����kI�/�9/>��GEV;�B�r˺�N �,=G�>_��X�2R�TIHD%�bMc,���¢�`j%�#/"p��x��[�9�@������e���~���F �4�m�ݴ}��\�v+!�:�:�6Ё�"(�( ��|�a0r��O�?f��G~m |7ρ_| �DK1��+Р�H~����Q�N�l��B���6�����x歗���o�Λ��~*�m�إ,Q Բ6�U�0�L���f�&��u0���Q}��+!����B���0�-0(��m	phJ�S���ǥ^Ż�=��ߔ>���)�R���0�X�V.�nT���O�U_��c`����Y��+��R���;~�6�4o������U��͛x����O�����K/=��_z���,^�.>��c�����؇�����=�#�
�J�S�]ip���U�����Ğ׮��}����k<��3H�.���]������=ߔiG,L�#0�2�ߍg�}��n��R����a����������#���n�}=��#��I� �� �"���tv��K�1"l��)�!�&��2�E@ �Ďړ�Qv,ᶔ�4<龍��'B(���������y��܏ZA�R�ع	Zܯ�,�F�>��>��9��@�߫����Hqυ@�H`S Sw�l?��ߪ�G���x��Щ@f�h�)���& ,P+@�� Y�+�W	�}X��x��/��_K���J��08L�?���� ��!��}H�@-���rK�&�\�2��HgP��v
|
t��&絛焥H�E;׫ԭ�jt�Ű�hv�B{�z��Z�d��e]�S�#�]I��OP�m��N����L�%��m�N�I�8���ǋp�^{3�ڗ�I�|��1���ԾdL�$D-�1�5�K"���͗���?�I?�˟���3�X��s�B0��91?vY|sV`RY$��WaL�2����0O�E��d�,�D�@?T�f��#�L��܉0�5	�S&@��
Zv�nm[3hO0��R��k�	0o�1�0�2��h��f�Z��;Y�����Z�t�5��B��=c,F�F���l[h͵��<;�g��s&(�gL�_�|l-KDEO%�^>�uy�0�4�á1Jc��a�M3h�kA�l$4��1Θ�1�M`�����᎖���а҅�h=.c�vN�c��:Sx\n��ao��nVF�z�@���\� gh�����(hL���T+ֹ�I�\G�&����t����/����������.S"bR�,���a<~k�	ؒ���\�w?��_{�s7`�\gح�!�@o��}�!�`3N<sO��<��{��e0��� '����JO�O��2w�-���ip^3��am�)QزRW �9�ۑw��p���׮�b�T+T�M
|F*	�y�@�Z�狀�x;:պ���8��B �rkW�t���Ƶ'cS���@h�mIVE�n%��s-�R 3�i#��.�ٶ�@*P��j'�>о��FS��s�K�Z<���]�+	���!�І�PIB�t�뜡�u���2�$�o���iڡ|Ż�v�O�*�Ϛ��JPU2"�ܴ�@��ԩ��mp�S��2���)�
���qV�mDõ.t=5��[���ҁ���J[�$��S�(e�$R���TI�Z2	��RJ""	�M�!TvgA�4�~�2���6Ԟm���U���ExA8���br�=\f��a���f�ѓ�0�E����l�1S�a=�c)�i�񴀭�(�z[���
6>��=
֞��0���!L&@��0������*,O]�,�h=�Q�c�9[��}���q�uK�2�F	�Y�T ���o�0\�m9J�8ND�ɧ�ć%�d9)Uud* K��R���ږxb�!�T|����]�ʋ-㔊G9I�؆� �^x�2����ro3��*���ע#S���-�kKQ 4� *��6Bh�`6��tBl�@����@Sz��ٗ�^��R�J��+�h�т�[h������\����M�����' *�� |Jn���h�҇���J�Ɠ�h=�{n��V ��D��[s�
�+Q"zq;
�V��j�}�,��TO���S�-T�qQ�r��P*-A:��������a�,�B�p�Xa��h8�#�h<ycڢ��%m�x��q��Wѵ� 6�b��mH"p�8����Vք���N)D|Q�뻑S�ս�P��0��{�_�m���Ǳ��a9\�`;����Rہ��rDdV 2�I��Ȩ#�V� ���t���g��]»_����G����x��;8q�,��9���n�O>ĵ'G-���
�9Y������n9z���YihiFyu%�S���L����g/��@r�2�N؈ʎ��us��zz����c��{���N4(�
_h�Q|�/,��A�*}@d�g��ɔ�_
`*ît��*Ɇ��jH�eeP� �R��i|��ǲ2�f�J*����E���� ҷS<�3s� �A����@)}ӗ(�O�HBteL���q���#H
�����W �?�N���}ď� ���@��6�Sc^fr_Kx�++� ���q;�!j����;sB�s��}���p���H��V��OH\˜ ��&`nWdV��5k��"}B�������Z(R���@h�x0�3N4 �J�#��
g�~o��;|M�����Q��@���1�\]�!�z c���R��g�Z�w�R��h\��E�<ZtG��vg��[���?�O>}���8�ݻ�^��k�O�ҭx�{��__��'w�s�A�����c&�e�Ons�?�_ɗ�!�y웰�/�޾����=��?���w�( �NP�Զ�{by<aI����?�w����y{4������^_��~�[�Y	+	i�X�@������ ��0��_ڜ�/­5r�n�E�6@�9H�"���JNR	>������c���*I��n�aSv�S֍v'sK��!e�/�L�=IЗ�#$p*�3r� �/^6���p��A�m2-��I(1@ ����P�x4v��b�i����RY������A�oX�zN�x}Ļ�$�y�.��_ T���V ����T����J��~R&�]5OJٗ��J�0��S T���S�7��m5	���+5����>@G:Gt�l�Q�QK"0S��V|N�&bTL t����=�J�l׽Y�>Z�Åpۓ��Lٛ�>����g�e�6L&|z�I�t&w'��}3ώ���g�7/5�vཟ?�����,�Nv!89�ｅ����u^���������ظ�����K]�AQ#�z+�)�R5f��	P�PN����X%!�@7�IX1Z�	|##G�mA�iC�X��#ah��1����X=Xp;V�ְ ��z>=Gc���e	MB��[��'@������N�U��V~������Q����U�P�����Z����<dV棰��;�Q�ۂ�A~s��]��;�;�B���8z�<��Ĝ5A��g���/=���k��`���j��ہ�	1��j�Q��r��=σ���4L�|YZP��0&����CǕj�I���3�s���������f0q���'6G�p�(og�6���.((������[w�ċװ6s��)���6��Оm�@(x�n��4� �n�݊	=�;�pL���Nt��-�
S�م�P��zo\/�>��U��&t���f/r��6)!�+��2~�$����I\І8DI��FB��C *^O%��|F�4�w��� �Ld ���'�ؖa'�w�)*õĵo�&j��@#��Z�6�7ukw��T�]�$_�"�F+ F h$������,�T���U
��74�8��A�m]�J�U�QI��dD��HBoL�'����h9��"��z7�݌jj��FT�iP�w�i�h�劣���C���H�+e�T6�$���aA%e0�W���Jh��
e��e�K�<�Ʈ|~��o��	:��у����v2���	�1ʖi��Qv��鱜7���&,'�a������g�}m�<��3l���z�h���`��ip�g�k�C;�do�Ԑj�������*O�,CӔ+��2%��"U� ��R���>�����M=���_���/R��G�m)��T�U��~��I�����ɽ���U캺5�ZQH��Q �mg��r�>>#P�xC���
��g�V�� �˦�
|�>I`d)�OiS��lD�@�P�
�M:��m�҃���h��ö^4��A�)���������W����>]ɇ����R�H�y@�a�9j�6U���Q�P�/�)�Z�|��G�R*�6	FY|@��V���N�>3��}E��Ǘ�%lf��#�S�x�+�Ӗ�!`�"d֔�yw/Z�`Kz.r����9������w�DEs/VD�c���_��y5HȯGrq��{�PڊȌ2$��@�(�u��\���pq%;� �����x�4�>y�o�������՛���+x���p�ɧp��c���Sx��q��i���a���@᲼��M�hڱeu�(��BYu��[��ߏ�ޝh��Gе�'����Ӈ�{l7:�u�����Iˌ����<c�N5b�KG�r��7v�>iE��zTI�O���˵�T����@!_�2K��� * Yr�/�S*o�:�УBp���[e��/��h ���Q-��<T��ū(�(t�o t�b뗵\�V��I�BJ�>��G+Ypm|mU j���h�l�hx�Z7�cg�?a������~.�q	�JPP	Í��@d�V�n�M����B׹���=���;x�է��:fK�`7��`V��P�<�'�T�f�7��d� m$���E �F �P\~Ԭz�0�+���T���B����I�d�����o]�&�ka�Gm��έ0h��U�f�]��4>g�v�$�o@PG�؂QUk��;G�.��_�w߼�7^��g^���_�Av�=Ww��'�p�'Qy��ht$ �p<f)^;B��`2iP;�N�$���R�jO��o�>�����?���2x����V�r�g-LV�4�@�j"������[����[%	Q��vx���UM,�d����ߤ�~
��X�����Ymhdo,4V�J��&����HB�����-���ݻ�`� #B�1�ӄ!�O��IT����ܣ�O�G�GI`Gk���GPBG�4�. :��'`J��'��AU�g6�����υ�)u��x��[٦n��TЩ ���rz�L?B_�*�`lx�=nҮ9@�T��(�PUx�xTyn���W��̺��}=����:�:������>�j��W���0��_(�� :� �I �LԒ̜�t4�1�o����f0H׃9p�O��&pf�co�.�׾\Lܙ��(	�Ǧ�J���$L�5T�36���d¨k�L��
wB�׎x�KcPM }���x����g�ػaɫ�<����Ř��NQޘJ�1�30�0�63����� �Z��0?LZ��%��b:ܗ�`�boL��{�x�c��	p ��y��n����������10e,L����N#�Þ���2�'��O[����%�P�6������%n0�?Q���,�����>��̄_�|�߸�)��ͭH-OFv]�zjq��[�=~Ɵ�7�Q)����+�~�Ǐ��?���a��J.����w|���(o�s���+N?vQ�����>��?q��5���"��%�H��qO8��L@H�:F�@`�
l��@j]>�Rb᷊0W�N��8�5}Mh?؋����Wp��M��:�\:���r$W墠����p��Y���x��+x��8��I�%F@���L[-t!��`$>8k=�>}�|�
�x�.J�1~��`��U>�Y�� ���y���f@����2��f!�#MW:�ܟ�5�Z���!��D�jJ�oeIBM�ϧ@�H��V$a�J�E�Q�b+��ܗC�:��0��gs~����-��)M�FB� �:	�� & ��z;�����M*���)u��<YF���*�|f)Yp#�>�2�iV��`Uݺ� ѶAP�̲��(��%�)�˔l�'	0'K�CJBl�ϧ��R�u(�)��$W�U��/ ��D-�U {_1���>�/�M�Pq���jPxd�Җ��P�JO�f.Q�	�nۓ��������Z�v���eJg*�/��ʩ���c=�
��F0�Ճ��!���c��XH��A[_���a`2B����/uM�Z-�`!�Ǥ���Fۙc��%�O[���{b"���O��t'8��`�3��Ma�J��2��JW��AFW
�O֠�bj�5��p��m�@�#ATB�%I���&��W��B��G��H����,# )�����%@��vU���|u[.A8�h�Su,�{�x��pO!�>�^����{QK -�U�h ��Bb!t@��2X�x$�JnV*
��Q�3ݻ�Qs�ps�Eϖ'	�j�P���*h��=�~�?��CІ�;�,��g��B��ى���p�ݛ8��a@�Zu����>�/� ���Cq�:�e#�`�RϧJ��@hU@`�,�dY� �z���C�A4��L�H�{�T�{����ǵ��	��A��\:��#�,{/�@{�.��;L�ۋ�6��Cg��]ڈ��1/h-b��a��<�\����R���|�L�Cla5��;����;�}p��{�O���w�{
=g.a���z�]|�׿�+���?ǳo��37o�g�A�w� !3ۛ�еkJ�x�:v`����ܫ�oح(���յhD��C8z�"��|����?���A��dw!�.�k�������y���E�^��ݨ�ڂ�uʸ�e�x���T�P�"���2,;Y��S���5JH��� �$�T�x���m����zy5��'�ECЇtVa���O؜)�I �)^PQ�2�H[��sC���t;%W�P@S�?PT�P�|�����M�73	o�� tAv��K��R���8��TBp��ᝲ#���s�bt@�~�>��s��񫈯̈́�'����9Ԙ�_��U0����U�è�u	��T�� �%ԢC2�n�8�o ޽y�OFxo%N��<>�A������O"�:	c��a��P�:�F����l� ���9���8B�����J�ժn-	��~������x���н����q���F~�5o�\B�w�zx�����Nc�e7E�ڍ�qٗ��pޕ��;1�5�wN��O�ᅷ��a�r����"
N���C��4�%	��5�
�]I�o���߽��	�7߽͏u�*�aBc,�vlR��T$�a7T�4:ݱ��HB�2,ƐdZK�t��3$�K�RI&�4	�#	D#�-B�6�G����B�!��Т��!^���I��&�H?�GI��O�&��;���xޤN��Q��H�,KU@H�_$�%k�L�V TD.C��G�~5�)Å�<=8t���oD��5��)���ۥMS�����5|�_T�#�)�)�p��T�7	�J�aP�>Z|n�)]B�@���^O���:Wr���x>���5��퍓�{�0i6��,>3��L���{�W�s?�u��i���(�:��I���ԗ��;6õ{��%Ϛ�t2�?�[�FM�!�ܱ	���Ncٯ,�g��ܧ������+��S;Q�[�Γ�4t�y���ki��s���6A���s��'���	/�֜��/]�+�O�sG?��S=��ߌҖ\���(ʌFx�
~ké������hlLY�I|'��:���<e�(.+��a~�����+�13"��s05, S�����Y����!3�5�[�cYF8V��`Cy<kR��=	%	H*KDZU���Ѳ�{����Gq����yO<ww^|�O�CvA*�
�p��Q<��5�z�*��8����X�%;�v��?~����Ox��-�7W�;���ן�����p�x�ջ���=���g��/?�������^��=��ջ���s8��\�sw�yI�Y/P�����ｂ�޸�@��l�3�W��>������O�le���|��O���o��w�Í�"6g#���~�L�#�ma<�	Mx����go��k� ��
��N�Ѽ�0���ӡ����+��>�0,���c]�2�d���0kk7��H�� o܀B�hU���%��Wh�x=U��P��/�@*�)��$4W���v+�@4��x@	����L��ߑ�-]�ʰ)* �6��F.���oA��'%uiW+�31,�m�'��B��^O�������[c��74�x@k�����6��J2K:�4�p��唡X*h��H&�K���
tF
Ӯ:D۞�
��K��tBf��bBW:o���W����h�څ�UJ{�n�� �$� %�Oej� A�����Z٣�g���@;���c=��a�d�Q�F0M{�H��0�=���4a��#]����PF�όi��>3��f@��Z9��XFf0�4��3��6��X3��'����p�����qJX��$-��4���	X��)��h�ҁ�;{��������'��mKf�>P���AQ��>�����e���,/R��@�/}<e9���*XU����A�Ųo�2\�@J��������{�p��h9ڍ���G�����x@3�h��� ���F��z��)����������0��cPBh�}@�/�d[7Nw)}@[Nv���\�q$�V��F�YJ<h�Ϣ!ϧ�h��2��P�'�70�3�`�"��3��PPu(.a��0* ���=Y��#�J?�M��zt?ه�[��ȓ�r
�ζ����`���Й��Q雐QUD�DCG?�jjGK� ����#�.n�Ƅ|�D���1�?�C���k�֢fm�"�����8�U����8};N�C������s�	T�GIg7�O��s�}��~�n�p{N�@Mg'�˫�Q%(nL@~e��S^���j\}�y|���q�O�����~�s／/#���-M8��-<�ћx������/�~��E�Ħ�d,��v��yJ����,�~��}mO�B��v��܁2�ҧ����,��l�Jg���/�b�d���D9��Us9�
p*z��>���X>��� ���3�>
@%�WdS,���`Aa0B���_������A
tJ)Yogf��2��������(I���0�0�"{@���<��Ȁ :q4"�aɶ`̉_�[@��IUe�]D�]V�` �xA%�-��kL�]���'�����/?���!�1��'�<nL�����/jR��HT��`{�k�(�A ��V��j߄ф�Q��vg"lwe©?;��V���p��;J�w~��?~��
�:6�(�`D�aX\�����~�$ѐY�zX�lUB���2N����%�n��~/~~?����Qґ�EY��[��܆o�Zxs;���ٽS���HC�F�;�s�~�,�v}۔\�����q�E�}���q���i�4��<
[�P7~��ԊPf޵����!�������>���|GP�<fˎ0&�*$����u�߯O��% �PZP%C���y�"�i.D:��tEݛ�T�J�"�6�Q�%��l��Q��%ϧA��'�����O�C��"�j~�D��Zh��Щ�Ǡ�}
x
d* �%�#�IX���L������M��
,̥>����QRE���F(a�<<�F�	d�gT TBz�$ݑ�p���} �}�+a��-���� ��) �u�T���x;�����>�&� T����Y���pw��U���>�멁��yS�;�Y��Gڇ<�ky/�>퉃9�kn�~�f����;�ӹ7S�f�cW�3�4���Ec£/.���|���'b�$&�:�[�6��}
�`���p�đ���(����K�x����7B�_��%>��U�����/���y���ߦ���_>ď�~�*���.>��]|��o��go���h�׀�wN�/_����3o?�cWv�kw5��#%7�Y��_�ˍ��I1H�؀��ؖ�QQR�fE	Y�5}=6�Ga��H�ٸ
��W"t�j�lY�E�cV�B�.�������_M8���$���i!��-ƒ���]���>o=�'"����6~���P�T���Zt�mC׾vމ�=ؼ5
c��`3��E8sxΝ<��玠���%��/JG#a���x��3��w������}Ͻ~�D���x���q땻��ҳ���sx�0�ī����'p��%<���
x���K�p�nܹ�'_x�o_S����i#\�3�n���^�k���?��|������o���ć_��{��»���~��|�
�J0f�D��x�F�r��Wlk)��n��[/�򽧐�]�1�Aw�$���0ttC}�L ��J�:M�o7����Y�������yJH����b��a��^-���P���oh����T�	�
B� *�)p%�� �$��X�s�x<���#z?4�'��)��?�V��)��p�r��I�����U<������� hh�znw�+}@���͡]Lh��C��Ԓ�䃹H��]x�g��'�κ�"^P��	IKJ�h ��>�2���vx;Z�w��?���+��'�Px�9��M�X�����|�`�����#!���Qp���:���b��h��jsWS���К�h�	]�a�����p�G�HGƺ�L==����02�����&��d������@G��:�զ��v]=��@�Ѐ0j#C���r�1�XDm-`mo�)c��i'_k8���n���8S�=�� ����v�;o��r�2�c�Q���'�� ��<&]�x^Y>�yC����d��vN5�J)�:��~��T����
>V�\��W�|�ڎjz:�v������U\�ChC^w94�7 *������G}@S�R�ܢ�L���s�
�/Ԣ�&�?����<ގ����PO�]oE�T@+�סH�	
<x��ڳ��;ӈ����4�W�x@	�	�v�����]�;��y�h:C0e��� N�;��ۻQq�
���p��7!����^rN�A��SNq�)e�����H=��T	�}P���#Q	�%�J=��f�=��q��#|JVV�2_��*���ڄ���h�ځ�n������
�r���~�faƊ �_�՛#�\L���Gf��:~�.^���c��kEnq���a�>PW��g	�F&"c{2j�!*��G�`���u`?�<�$��.v�:����q��M<���8|�2�z�ѽ� v:����ap�q�t���%5Mؘ����zlJ�G|z���P\݃�Ǯ����Ş�p�ғ����8�ؓ���+ /@пj�TX��6��@e_3rZy��bKe"&��w�\~p� ���ys}�4v>5���h�ف���~���H���Y���O�%v��S@Q<��ҟ���j��ҳҧ���.�塓�g�B./�j`U��߄�&�Jǚ�XL �����>���ha�J, L.�Œ�p��)��K�kz�E�����
�8�����4N�	==-��hC�/2]C���	��6II�Ԃ���L5Y��]�I��%XL����)1'c)��Q˱P��In��q�6�Hf�������@BK6N=	Ͼ�^��E<�֓�h��)0�0f�aD�6*$|���Ii(��	��'�*�~F\%�P��ÆhX�l�}�68�h�N̀;_��yp&�ϭM�W�Ɵ��?|�Wi��贈�١*��є �e�f��¶?	�i�Z�$|v���}�0�6v4�(ۦuXؓ������7oỿ|���}y{����2��9�}=�r}��$��<Ҕ~hN4�'�IŤCY�!x��I���t8Ȥ�]�Y}Yٙ�C4X����S<��+��v§".4h�[�,w�a��t��y�x�o����k~�g?���5�W�)4ƶ��#}@w�B�3:�Q�VW��GB�%#KS�� 4�F>(���&���t	.z�[	��x���_�6��	���R���-�'���5�0�E���x2n�t$�S���M)	2��dZ���O$�p4�#�K\�W���Ա<g#ڣ���zG4!XB�`y�XW����aW]\�3� ��������O���\F�̄=S@V�&ϲ���TY^	�%�@G5	��%�ʾĳ�R-i����a�^�� ��C���.�yl�{y.)ɜ;l�@,۹��=[0��S2�r�#�/ٟ7�EiK]�r�4��6i��>5��<.��<#������s��k�� �[�y�����<��T���;�����HM�M�%�6���ga�`
!4>����to�D>Ǔ���sNOڱ�v�a��i|V&�%q�4L�2�|�Z�<6n�K�:��E�ͽx����C_S����x?����O�������&^z�,��ww_��;w��'�����8|�͇P�]���U�;�;��a�DZ��#�`r)��.���K�f]�b	��1K�u[����ik�9ᛂ	�˱<rC��8jV�cv!�?v�s��0� �ᇩ�P�Έ]� ~goZ�����2%�kW����|��V"��i|OW�A��.�q g�;��=�c7� <~54L5��G���Ko��o<M�{����V����9u��ĆmQ�s�w�zG�Ɖ���ڗ���O^Ɖ�O�����i?v�ۍ���>J��@^ڇ���+��>��?N>փ�����#8z�^ݏ���n�N��v����^칸�gz1@�0��W���q��8r�867��j�;tL$HN��B7��#���^��/���ǯ#�����`�됹0	��2�����>�����;~	<7-�Ǻ�������!(?������#	e�j�!��'^ϐ��C�UE�S�E��T`S@��0�J%$J}�!��:��	��I� ٶMP��-��H�C*�����$$�@4q\O������;���y���:�V�rM���҆��[6*��TiX��4��ZM�8�a��� dFJ�-ʶ��E�l_Ӷ	m빝M�ߛ�$z�.e�g(��Ѓ�|�L"��,�I���d��ҳ5��Py�Q�B�h�SBis�}_�b��E2�
m���2�
jh:�P�R��P����xq/��}�^:��K�(>X���	O�*�@���V���2Km�"��x>3h����J���EBk$,��,XO��({cY�B�\Z&�1�p5Z�����cD�PFF�����	�ff&026����2=���fF�AJc}����i��DٮM�MK�ۧ�t�eB�� ؎1��8s�������<'b�tgL�9��u�=�#|��y��Z��$yR�/c�*QP&�;{%P�a�i��x����&�ϣ=�)!���夔�#�GH6=,u{.6���n/>]��3�(!Ԧ�:liۊ����� ��Fá6��mEI�#[�ұ�:kk�ל�-��,H_�4$^��Q*m�4�fa4c���<Ng!}g�v�a�v��m�FŹjf#ڞ�T�`i�!����vE* mU TDU���E��gYs�a@�sM
�6�m}$��	����(?,{���WOc�S���7��N�]iE٥:�XF���S�e�O�%u�J9_�������� *C�H]�q$� 2J���
���A�z�b����a��҂���a���ї�)a^�����,Gx.���boL[��������9| Ͻ����x���H�+DЪp��cϾ�(�l�X�m�@��+h8����x�oh��>�������h��Azq��Q�Eh��A��n�=rm݃h�Ğ�p��5���{x�����_��W?�����g��� ������o����R�^T���~Դu�}`/�=�sO�����h�׋��Z$Ugbm�&�H
�g�,,J���O�|<{�������t�� ZK �K� ZB -:���� =��E�F�4(K��@k��v���<U�Y��� ���nۓ�(����B`~��Z���J����`,�Y�Ey� U�z>�C*`*C�H��@.U����p�;) �c0|Y�C���2��>_j,U/E-ֵ���򄊇TCo8�����1?u5f&/Ǭ�Ř���ǷB�bkpy$�jc���%����T*ɋ�捂�
\y�n�xw�=�ۯ\EN;4��1�O3����m��n\#�A԰,F+ê��,uQ0���A�:���;��ГWI�C ��} ���+ǜ�m���e|L{���[���W���p�^;;���	;a�-!��0�;�;�`A�����D8$bB'�k�؞���/❿~�/��%���n�_Y�;�1��3�7^�|�M�K�� ޝ�����g|�,8�Cl7��އ�/!]�x�����x�����g�Pt��c0�1�F4�U��v�¾��w$��(.��Q��^<��7��������d����ԦMϏ�)�{]%	Q,�����-B��$�&�7"0�|H
�
,=���(e�F¡
FU@*P���$q�fhlV��a"���ţ&a�2�x׆BbEJ8l�:eȎ���-R�r;��e��yH������܌$\���0�b�J܇�����,+�c�
�d]B���(Ϗԕmr�a<��y.���x�2��pB�0�� /%���s*�*"�J���x/��D��c�������$�G�  r� �2|�#|�c+�(PK)u5��/y]�/�/����s�#x>�G�|��y�R���<#�y^�˹�s�s�>�Z�k��p˞͘З ��DB�{�ʛ�1���}*���Qw��'�/����w���'.�[0���
�g>/��֝�
I>��6��p�qmKp�� ��X̬ڄ�+=x�����w/���n��w���W��闎��K�q��.�xbv_hD����N��A�j���5�%(��Ƕ����CJS��Q�K;������@7L�s�;x�t��,7�ΞO�I��
����o������e�)�\��nΘ�96�m�����0n�3��s��gE�NĸE.JP���p����9�5Qs����`iJ8�K�`s]Bc^��Z���Iۣ�Ń��9؄����򃑫)�Va���w��;�y��g��@�{��X�
���0w���d�����|7,ٴa�O_�5�шʊAdFV�"~%�V"�p#6��پts�Wa��`,�K�c!�{N�<, L�b�K��Y��,=C�c�rO�.�
��S����`�������~D���@�t��
���
�`?4\;�w��3�oVo#������1~4�l��b�R��>�m�(�&,��5r:<bf��,�'��bkO"�@%�� (��
�6� T�1C!���Ϥ2F'�U<�"ip��n$Dn$��X��dH<��T�q�� �
�nݑ��g�U�����mO(�S�t�T��Ghx+���I���Ff}VׯU$�ƶ������^��窺�-�������8l۟���eJ�G�m" �}�Dɉ���D
��C&m��e
x�@�@ehł��(8R�on%���"�ȸ�Ŵ�
��@�	�JR��CE�'4�\jB�ӽ8���|n��`+!���_��Q)"xJho��2�S���{=E<��.�G�%��=(�>C�����~ca�s�w���FB�hF���1ц�	!�0�k�]c��~#cS#���(�!�Ӕu+k+x�x`q�"̜;';��q���F�!��X��Z
�겮7�+�W`TF&�ܶ,�X`��5l��bj�<�15�	n�pY���u�XC&�/��O&���M�%� ��ذed^'BgmZ����<�J�P�3XO'�* :���.��=��PI�Tx�U��P!����6��{�s�=���u�O��t�!����,��I��ꭈkJ�Vh���C ���l��K��Ȥr�Q:X�ʞb�Jd��z%��V����Q{�=�L	��� z� ������b�.֪ �,a��֣ 4�`)��%�)e&A3}PFU�IPa�Zj �z.!T���	�tǓ;q�8��$u��#��3&�a�3���b�"/x/����A�Lڄ��8p�$���G|��?���k(��AS['9��g.�e�Vu�����/�~� ���g�@ }��p��cx���p�γ�yh/Z��Q�T�ڮv�:��C�	�M8p������\O�W�/�W?��>���<p�~���p�Ϋh�ݏ�v�0N]���7p��y�r矾��S��L��DTNlƌ5�����_8�C��B��}��ͨ�M[}����Q}���^�������&}8	�j��&$J�+	�8��L��2���W� �T੆�JE��n�O��y����%����v�s��W�Y+1?{�#T-��e�T<���C]��Yq�1l�Hh�h�eH�����?ij�O�42&�i���@F�|9Pu���0�8��s��9����sa�J,)Z�xi����V�nb������t��7͆��5�'���'O�֋��ĳq��+(�.���n0���Q�`��k���Q}J�@��W�
��0��Au�k"����b�Lm� �έ�ۑ�Iip�K�T~��3�iPnŉ�o�K��O������n\J��ď�������efGp����a�l�Lm�8��4^]v�ÅF�aնq���Kx���㫿��}r���1�l\�`b�:��n�GG<����.�o
&��±#n,��ʂ��lL�����'si0,kLB�C��իx��q㝧Q���	�ᐴx��-�Q�
�������C~"vW���8�������C��6�7�p�1�o� s�!A���x>�"�r�@V��-\�B�F;U)5��E��7�C��P*",�&�R`��#0*�?�(M���%����IH�F�x2ܸ���r_zT]	�~�	�Z��vݯ���D�	�Z������h��0�G�}$�Er^��'\��˄ŁdB+��5R��9��J<o<V�.�{���������o��o`��y��  / :\~����Q@���k�H@S �`(0��Rr�&AQk�P�!B��@�x�)鯫5@�W���t.Yj��?���̻?���}��F���{��D��r^���~��&u}�R.���$�"Yuo�asҮ4��J�S�FU��
|N��|zj���{�M�;ՉƮ]�:B�&�6'v�)P�ڵ��<��j��hL���w�:,kM�Z>���%�{uE�b�H]�e9��(c>�$�"h�a�F?l�����+p��� �����5�	S1i���t���,��j3C����b�̬u`2FW%k�,Ńbnk�	�д�x�l0n�X�r�����M`�a�iV1�#<,��e	-�1Н>�~�0r�t	[��aL(5����vЛe�9�\�
�oL������.p�}�'l��c�BL��I�X��َ��6�"��v�&+m~60��Q���_�B���i�����n�����l ~���3�F^�0�a�Q3���g,FN�����Hb �5��r5��ɦ�n��s3����Jv���Mh�k�밮��V�v#خ���9s���8����z�U��y�y�����k���ӷ���)��7#�~;³�a~|4�%�`a�Z���`L��߸E��0_I@�=���}�ئl�LQ��T)��~���ʈFB��|+��J�[��Q�G���I]��m��q�)*���e�OQ�|��~�,Cp*ueXPY�����:ex���H��5����Q ֲA�@C	��'��)R@T�%���W͓v����c#���
d
|���~�Ei7]�$�*I:��~�@��M���E{Jt�0z��Pt���R`S<��
xB��)ФR�/�����!@���LP*8@��&}I��f?Q���ۑr�Ʉέ{(\��B��l#�ύ�}�FO6���ᱴ��4GB��x<����@3}��#T꙰$l����~� 5�!���c'X���aQ�T�V-GDL8B�W*@�0�~F�ϪTKW�����U<���gT`Ԑ jJ5�2�xgsL���is]��g�}�$�Ϟ�)!������ƍHHG����u���=Q���tP��R�����Lݗ� ����y?E��Z���4�׷�l'����Jޙ��=h�Ё�z�}n@ɂ��U���$��bc]��&�W ��'��JP���ܖ�z�|�M��) *c��7 Z}�5�B)�ڄ�3�%��v{�ه�����<�ᒄ�֠H�%̨�( �|X�Rf@UAi���%��(���ԏ���#���k�8��	����­Ka�;��`�B�X ��3�2�"�!"!�}m�����������ֳOc`�n�<w�����~�w�F���4��̭����+8u	�.>������S��ʳO��ŗ�o}�1N]�����,.Bk�N���W��S��O����[Ͽ��w���×���<}�-���g�����w�Ko���w_ĳo���7�ێ�N� �<a�\����4�b��&z�$��t�O���z��l���MՕT^���+�t�ż^��,��'&5|f��'! ���ڻ)��@��O�E���n��ٲKVbN�R�#���#tB���U�t~N�#T��~���:�0+J�bN�R��rĨI4$�=AT�/F=c(_FzF�J�#���Dz�@��1�3gk��,Jü�U
���vyi8���bEy$��֫>j�C!�-[1=n.FN6�O�L�����ϟ�շn�州@�Jx�����������\
��e���n�
�D�oh�*�U�B�2z���k��Ic,�a͏���M
�N�O���D�4o�y�Rx�n����Ň����S<����8?�����*�¸�Up���X�	c	�&���ph�A#a�%-�A�j����ҭ7.=�p�ᰤ� ��|������{���ʃ]ٞߜXx䮇k�LH��G�fLk���eX��+c1���6{5�rC1��>=阽� �� �|��|��|�"���8���@di<�łҍ,݄�e�XV����b��y��?|���xo�.���}ԟ����P8��`l�
@��cG0�%	���Ft���V�V�j�S�݇�_kX�o�!�
��:� "B��0UI�	];�Wˑ�2�>B�r����-c�n��D��s����h����}�k�V'���a������� 9��祙�^�aД:�	Hi�J5����9�X6,xM��5\����R����8o����	Y���0=�N��2�O� '���/���!�*��R���(!���I~d���%��$R�~��[��gt�'AK�z�J:��	%\J�OI>4��c�����1p�r܇����T����3�9��o�Z���-���LHO^_m9^�gx�4�x����@�_����z ��0�`���2�ʾLL!p��P����/QU���[�D�2���u�Q��rڑ��6>���f�Q�i�R�ם���M�2X&΄�FOFN��j{�:�,b"�W;�$�	��Yr^�WN�E�4��y�d�4�x(�~,w��"g.��yN���TK�Y@�������}¦�h=EzV��5�.AT� �=Z�RG��&Σ`�6n��Okx�����m�����~�E�Ӝ9s�S�T
����!�g��sl0���𹄽@[�,s��90"`,������V������0���੘���TMB�p�����},1��F�\]�c��X/��E.\~2��a���v�qjx��0�1���J��,{�R�y��g��0��J}$aY'��x��N����<��<��`��6Wq?��y�Y�-pT����=��s�0r�x�-rĸPOX�{�8�:An���1 \�/� �{#��G�����ǉK�q������+������o?��|�����m\z�IT�m����������a�ڹ�[7��bi�jD�l�ZB����O	G�U�(4�ߝJ�`��[5�JX�tc���T 4� �LT R�b@72%!Q!S��mQBm9���OT�+* �)������wZ	�%tJ���u;8M�tmCT����-�F��)�)�)�O)%W`�A���/��3���� ��! ������T��"�J~ɉ"6s��K��r�I�r���=ۈ�m(=Q�R��^����g��$0	�Jn>����Hٕ���ٜ.������8�(%����m%q)���y5�u(a��uq����X޿&��0�cs�Q�``�}B��z043��S�6���1یahj#3�Z��F���Q�q�����	��~�1k:�,�����<d��X�K`F�t�Nq��#�x�%��}6�[��@�
L�CJ{��l1�6.������S1}�4x��������ڵ�۝�2y�x��ߦ �r>�/h:�3�@�r���[x��T����S-u�� ��������Oۗ�ľT���!�?�w��J?ZN�@�j_�g���B�5�!���M��
@3v�`�
@�v�����W땬��+�o T�Ɠ@������{v?�E��]g�Py�e��Pt�h<�	5�Ђ_��Z���:��J=S��G���J9��<I�a=��J�V����fBסW���g�|�A��`��)?�N�n�i�\6�0:3W������ˎG��><���x����_����揸t�)t��GS�.���|��EׁS��?�ֽ'�0x����<�o|�	��ᝯ���˗нo��?���y���;�}�?	�.?��?��}�A�K\������'/�o�A�y�E�]�-�����+�`�pG*R��A�a��a9oGbSZ����q���h�Ս�uךQqQ�����:_�kE@�X�������~�O�3�0����7�����M%�j ���D���LD�o�Bּ� ,,$t����pGbiA8�>@%�V T�p��-�F�¸|8VD!<7aIa�Z0����2�T@TCK��!�\FRc#=����Ѐ�t@���|�5���b� c5f�/�bcPY���%��|�*�C�U���0�!3�F���?���{|���x��ǔp�yIK19q>L7�a$!td�h��,�~�s@�^P��Ъp��F��&���ٶm��Ió'�}ɰk�ǆM0&<�D���x�w���µ�7p��q�n���u�۲�s"1�u��L)��!oZA�2b0���-;.yј@��-��Զ$�иX֞���/Ὗ>Ƿ?~��߻��#}h9և�0��e�=}E�waCo5�������ۇܓ](=ߏԃ�Xڔ�9-)XЗ����Xޚ��{���_?�k߼�g�}O�q�^{��}
���u���O��_��G����%ަ���x��Ɨo�?�����v��0�Ց�j���x@	,��k�ߵZ�)��HJ��x�֐��a�a�Wj��_WC��U���R�� T�&a�T�:�4��$A0� K�i�]c��>��݉�h�~Z�z�=�f�4�f�������@���hևAc�
h5�È���}j6�?B"aT�F���phbF�>�V��vSt[b�߶<�R�6��htn�^�Fh�]�f�:���i�تJFD��$�)c{DҏR<�q���U�`�?���d���>��n��N��)�]��/mcw�b5ao��g��0fJ(S������b0I�7������m4�o�����)�L�x��L�۟��4'�b���M�1�?�����m���ce��Xvo�=�Ł 9� 9��"@�ߙ ��Lٛ?�siL.���d%�(\����K9��e��\���c�`&��b��|�ܓ��4b󽼀������>�?�s�)�R��O�:�\�9,��mTB��W�b�ܥ��^��%����Yw�c=�C�~X�mK����
�����y	̣g�8�kf`lL �F��j�'F-r��w��C�1�v4���Ll�a4��i|:.�̡oc
��4ZY7r����9XN�)c��9��F ���-4g�f;@k�#4����-�ǰ�l_>#�MĈ�Δ�"Mj���Cw���M"DKI^0�o��RZEx�H�!S���p�;�|*L	�.�K1%=�b`:�ް���Ʉ�?O��iC��˦(u�E��n�]*���*/E&a�0���մI����_���N��%�s�Ҙ�o�ʃ�&$G���+�@��E�$X����_����3���m΀有��uDB}1Nܾ��wn��5�'���ӏ�޻���Go��_���^��/^Å���{;į�o�%�S@�<�ٴ �y,�X�����*�����kU �ii%����j7 �>N	�U��
��O����ئ �|k7�.���]����R���A���eۆvn��$_CL+�C�%x��NBlO2�**��G����Q�4�&0J��T@�N����̣B�|d�zDwmB¾t��@�x=e�BBo��>��C�������'*Q~����*T]��~u�N6@i��� a��j�̒�6��L��*����2��$��!ew6R���������R�nI>$���\nG������Af��Pi)C�h�@H��4ѻ��*�42#PZX���
�ƌ���5��X�FcƎ&<��(+�Y�a��&؎��qp��
�^�𞢒�ez�|�h�r��	Ś�D����E����D�5#�	���UK�[��i�uaam{�q�
�� /x/s�4>�>��X�u6b�G!go>*N�����S���i�6��FiGx^�Ε>����� *@+	�� iw��}H�IG׵��6���=��ߊ��
|f��`Kst���{	ޅ(�/DM9��I�*	z��q{Z'>މƛ��m���B�} �E*y3	����L�lE#A��|��j �$D�$	Qϴ��tz��)!�{� ���Uכ -&�J���@�+)�	��P��Q ��OB	aR�J�K;���C��!T`S T��@�) *�I�(='�r*!}e�����������X_�.A|q�7��S�y�?|6f�BCfa�ňM]���tt�������������O|�����8x��Z{P�c����{��{�Qل��f�|7�O�ƱK�q��9��tן���W���{'�+���ӋϿ�?��p��c��߇��^����p?G��g�����w.�bg-�+3��$	��xKf�]��i�(�׀�/�Ǖ�oc�+���dj�4�^hD�Z^�r�g	�g
Pp��xO�&4�Z��S��S����)ա����X�l��B�
@�O�sJV\�7J �$G2N� ���9W�H+b}�`*�aI�j芡,�!Jh�ʲ(��C��(sW݇M>YJ]IJ��'e��4�`5�UDcyi4V󅹞_jc:�*��.��YGcj��Ih_�Ì4��
:�#���BMM�ol�x@G��E !EVSV`n�2%�V�>�8�.�O�n念R��5c��� p��Ѳ�o��|�6n�:���<,LZ��@Xl�V�<�L���E��Z
�� ��|���^	!�l5�x�t+VC�B�ŏ�}�V��#"}@m��1�e�6�$e	�W�ޏ�y�>{O�rW���3w.`��!t=v�O���3���k���x�������go������/����bہ&�笁G�&��D������2���w��G��'������k��P����/|��?�½'p��[x��{x�����?|����;|�?㭿~����Қ����݈���|�<>����)>��|�����?P?���2Fߟ��?){����ワ��so>Eо�sϟ��O"�@	&�܍��ikLz���M��>�P�mFv����X�]�P*�������ai�6��V
|*"�
�v�Uy��*�Q�}��w�6�z��X2��o�����]�ktz�0R��
l@5�ē�&q�S��8��G�G�؆�D�FÚ#0L�o"B�}ՇB�:êWA�<�=���1~��VE���3�{�����[��5p��;Sz�aK�і��}S�%t�Ӭ��!:���5��Q��a޸�o�x���̈́��|��C ��
���0��3ʂ���>�;����s?��`��L�D��3	�� ��uhڂ	5`_�	Nu�1���5X�;��ٞ
��4�ȇ��Ғ�Ȼ+~��ʼ������¼�����T ���#՘�m�v���Gk����ݙ\/���ǝY���H�gK"<��aZc<��Q�n��Y�ڭ�O���dLoJT��S��+�ӱ�)�%�����4>)���*�?�Z2��!k���%�}%ذ��=�XT������nV��cEK�7�r�4sZ�%IX��ɧZ��,�(�ƌ���^��L�X����D�������i�BL�[���uK\6aʶ�p���i�RL��e7aL����a�z�h�Yyc�rB��)0�����?��nca0��60��,�G շ][��Y@מ%�K �q-«ִq�C�a*��E$�j@�:*Щh�P���H}1�t�#�� �� *P�A���bF�p�f�D�u���-s�V��"=B�� ����
Wncۦ�<f:�"<�2�۟���F𝢔&�a>L"�12h*F��՗16Wr���j�6Eʰ'l�Y�=§.U�5	��KC§!�ӈ�iN8�L>	�������u�F�>����^0���ٺ�0	��� '�pF%m��~�
Ͽ}�n]���p��i�?{{�B�4ف�C��,Cx�:�_��s	��.�aYj��� �� ڸ� ��|�WVKHPU8n��h5����pٸE��C�����,��P\��
x�!r�r=t�x<�$xr:�u�)@+��n��eU�e�Qܞ��x@��CRBq��Q��� �J�@�T�|
T6�*	�$�V@4bH*��:U��!	�F��*I��e��@��e�{B�(�v ��e"iA�6X��:pj;���Py�	��i�_�A��F�T T���w����!C�HH(�R�%Q�xFs���>��$��6��}9]��*^�RB����E��N���mA��m�QSFAo�6���`h>���	S�����	���M	��:���3��'���v��st�������� ǉ�p�\�&���Y�P�~��0�m�����3����N��p��I.N��∉�1�c2:�D�c[r<�	��c'�Q<���S���T�S�#j(ú�i��s�L&��p�������43���{b�z?���#gwa��v+�P(Щ�M���������Ð�@�P���J��lnK������ݡ��������G�i�f��)H��@�.���F˩�hCVg)���+W��E�o����� 4M����]�H�����wf�)@�@��
Q�[��]5�>��/ժ<��%	Q+a�� JPT<�* ���Pu
`��A@kN�)�٠NBt� z��y� ;��t��v��* �@�l8�B��U<���ޫ�ٳ��Ј�kMJn�9>���ϧ(G�C^�G���[�x>��`� ��	�>�#��Yp�T)� *`Zp��g�Q|N�Ub���_nA�3{p��K8��5T�Ǭ�`<�c���g�t̍��L�����@,�Z��V !7�N��[ｍ?�M|����
�}��������g_���{h�}݇O���1�:v
�GO`�ɳ8E�<y�*�<�=���g��tu���7Lo7�}�e<��s�,.A�\�uWn?�s�]A�����X��1��6o�#0=r���`]�6�>����ɷ/a��C�}~��B3*/�(!��� -:�s��{�����%�>���+ =6~�+��*`�k���H��]�0-��/�)Q񂪇nϧ2��' ��>ZIB$ *�%ūT��J����#�x�R��>�> �~
�ʼ�o����s���HDѨ�X�4l�]���m�J8�v����f>� :��Cǈ/W��tLu1�XV��0o�2��c^v���JB�~�"��U1Jؐ|�⺓���\L
q�d�͹x��������cQ՞��c
�!}1�RB;�"��d,�N�2��B�J �'D閮�vi��W)óX����y�`ӹ֭1�B���e�!0��:����;���Gx�����o�w�?����(r�_������'�3��������`�?|�ᗯa���}m  ��IDATxJ��h~(�(����+_����?}��p����O��C��W��?⻿�7�~�߸�g�z���s��/����{k�s��� JhXNC|�+�~�O�D�/�� _��>�����x��7��o�_����o~�6~�����p���b)��W]$Ad�Zb`F83Ů-0O(Q<���S$���t+��!I��߈P��N>$	5U��>����d;!T��7j[��O�rD;�T ��h�'�-j��5$	��\�bp�Rj
�օA����H��0�fV�p©����UK�!x�	�����+`ҵ�'�؟���ᘐ��1>j6L#`�& .���J�4�+c6.Ĩ������u�`�~>�7/�M�j�e�Ö���	�����.��{s"|}S	w�4d�GaL^8�2V�2%��A�����:2H~�t��`|�"�nX��K06��Z�q�0����p\��Q0n�l��=�u�S��B_�:,-ن����NQ��Y��:LO��Ը����k�r&Ƭ���r���f`\H ��a�܇��q��Yp��mV��>d�/�Ũ�n0��#ʐ��e-��M���0��[8��u	an�L����{"̧9�t��RZz;�{����p^����.��K/{X�:c�LW������6+/E������N�w��Л��O���x�0���ct��4��=����}'�z�6��, ��KX�¸9^p\4SW/���=��^��u�Q~9�6s�b�'�4��3'��q�쭠oK�$|���Y���̡Ei���4
���ɄP�&t��	Иi�P����@�2�]���
�:`�s�'�\�xDG65��a�#�'tj�`�̓�i��]ϕ���ÃD���I�D�dE�aϑ!�J��㨙�$�j{�x\`�i�����9\g�J+�)�j>E��YQY_��By߇z����J]d��iG�R����0�>��ft)n�8���\a8M�w᳿��'_}g�����Ϣ�`/
Z�cSE��Ec�֕��%~|�d��5�1-�~1�J&�ŉ�6&�P<�k�7Z�+��be�!��O	͕����OPɄ�`\eh>9o�.	�$џ��@�\J_P��2-�i��'U�! =@¿|Jh�UBy�m�*CI�D�!V"��F��،� �R�]\�S�@�����T�xH�O�]�T���E�
��t�~	�%�߮�લ�f+��"�&0�mK����$!�W��\��N m�҅��MJ�B§:ۭ �x:8eZ`T$�G� M%�n�E ݝ��y�r�Ö���H�r�\�@Ao�-��;�O2����[j�Ђ2!�R�&�7�KFOsCB�)��-���q6�	�FWW��O���d���2��S�0��^��/O����z�5A�NP�iX�l�����~m�t�� {�ُ��dB�t/��y�/`:�ysY'[�m���:)�S	�5ԃ����������w�l��Z�}�3f,��9|����q�[�9{���x<sOoG� �����~~��S�S5l>��ƫΞ�1�����$�����BҮ$�LF�\���<܀�]���L<�Y��܁
�5�"�8�u[��#UЄ�$�	���s;��(C��]y,	���(�U�*n�C��>��P�}�����5�PQ>o�G�P\4�"�>@�� ��I�j	yۯ4(I�м�@�C'u�]b�������
|� �9��ܓ��'�qKQrV��5(?[��[;q�x�ۧq��)��'�k�/?ޣ0�o�,�@@�,̦�07t.���ܐ٘�*����M8{�4�|����?�(��+��������7_������������/��g���/�#>��;|������S�)���/�ɷ���W�Csws2���q�z�.Nݼ��v!�����L�Fpr(��c�ZEϕ�kQv�	�_��_?�co���ݽ�{~�;Qw�/����XEߎBy���L�f��h ���7�/�ľ�=�j����P�J��2�[�v5(�P��\��m�4�/��1�_��" ��@'�eWm�AHy��c~vff���M]�@�"�B%��Hh,�0AE�XQ��ya���8k�6"�3y����Ǧ��Y�K�t4�4��GF5��(5j�h��4#sR+}S�(��0%wUe���ZЄ��C9=�F'���K]QЖ��>~Q�o@ys��ͅW�x��$s�h�������+aPB�,]=B��U&�U0)è푰���E]��kEY�Ͳ����#�#�����K|A����?�O���W��O���?}�~�� �9>��#ޯ��/?�w_|�?}�%�F��G����ba�:L�_^�E4v�;���L8��[����㳯^�<���{o�u��>&�~������|�������5���x�����>Ľ��Dϭ�Xו��ɘQIc�==��]n��'/�֫7�����������t��z��!����<��^8�k�]ĥw�(kGt$��4�u+1�3�:�N�g=�wn��u[�-L���%�@I��~���� ��F��;����������ձ��G��$HJ�0��fh�x8��B$ˑQ�V�&���tD=a�`jF��LT�i6H[�o4��9LOJ���Q�#�B�Y���^L%��F� w�GzB{�$�ϞK_G�F4�GC�e��9p��:�n�7�F��;��8C��	z.]���h�;�y�l�7L��H�,VL�u�l�,���2_��5��z�|���h	�����a�&�O�g�L����~�'N���=�Mq���8�X�A{�	tƘ*�1�X�KbB1)���NG`x|�b��$X����g�2O�k�f�	�`�8�=]`�C��p���-,��x/W�M�+w�q�&��i��(���	S'b��3l�L���w��14�F�ZÂ�t+gX9M��I��uq���JX���=�]�0�Ɨ�h�X���zLY�k	k�q�@ck���k�1p��d��s��5�L���`1��(2���oe	}Sc�ӆ��t�,`8����Xu��<0����l�c
X8�c"�n�FDm\�е�X�*���ĤiS�8��M���d�Ou��[���9N>.��p���#��������S��0v�q�<	�z���$�jٙa$�����9FN����VО6Z>�1|����!�R�l1l��DG�!tε��@[�������$��X,�
��P�e*#L[A�6B'��`)�S�F(t'4WN��x 	uZ+�b�4�L$@NU$L�l_.�:Y)�M���Ea3�2B��t	�Z\V�C5�Qڴ	�#�q]J���*�yzܖ�j�Q���F�ψ*E��(�����SzQ�G��a���~�����7�ǉq��yT��b��PL\�x���M��l>�{���|y�iCM!�zG����9�E���D�ӰU�FJ_OI<�( ��7D�t@#k7"�f�kֳ���p*�� �7 +�I �@�z=T�7�H�Z�$:�l���X�-� )cy)�
o'ն	��,<cv�c]�6�ݑ������Jh�/��xA	��R�5|�b��x@7*�\@+0�Cc��BU�>���qX�m�b;���+���Ԭx@���3��ͨ:�<��$`)! �+@*9QX"��Br�-`s0){��H�+q_R�� ����^%.�a���-���=,��a0F��[�CS�D�%A�\&�0eD�4�x;��.s�;H s��<��M��d�TwL��}�dE�S���� �Kӽ��L��;�U�%.Θ=�!�!`�ڍW ���	�����^r�(���ӑ��S]��[X�)}AE
����\}I8i C��.�K&��6�1:�l��3�0{�/歙	?~��c|��ve�Qϫؾy�w��X�Htf����w ���C�� 4� �m����&#�?�g�Q{�M��Q{��=���T���ǆ��� *Yp�Z��� ZB �
�%�6<֌�':}��$]�d,��e S����W �'^9�]O�@e5x������	��ԙp��
:����Yp������ǳ�u"GѼ��Ӫ0]�U^l��ډ}�����n��_Bϕ~����l�������.����s0g�\�/���<O�Z�E!�_�miqh�j��+����w	�_�ϊ�o�?�:����/��Q���7I�������?�(?����	���S��ߏ�N�P:�^U�M��L߈U��y�	\����rd��-�i�u����e���~�v>����S	�m�.���	�(;�����Sr���������7���_�׀/��%���.zD��+�(=W}?W-�'T 4�q-��/S�	�..Z�����0��Vc~�J�I�?���镴 �)�r	�e��*��ץńϒH���AH�sziqr��Vae�Z$f�գ�p-6�%aΆŘ��+Mh@)C7��0�sVbAֲ� 4D��Pu?�����u&lVL��U(h�����ƛ�<�K����1��]˼�0��Q�rP��4/H�jP� �~�*薄`dI0�
������U�C�k1���YM�*�`Y@P,�F�SGp�������/_�s=�g�yw޸��_����_Ƶ����7q�yB�3�p��)�y�.<}O��.�w���k\��(L�^�I��+�8��M\x��ދ��;���>�1��W�s�;.����Gq���8��U}�4�?s;ߋ��P}m'���`1��	���Tl廪���3m�9X�d��V�����(?քm}�H�E*%}��h�̩����4Eí=�;"a�#B��R��(�n�����JhTI�#\\�aI���RBV��K����{��oBu��d���-1ٺ#��A�=V�N�&�I�T$�I�/�JhT+�{��bM����ZR�f>,L��S�S�r%4˃1\��
eZ�xFf-�F��}B�t[�,�B��y�����]
��y��( S΄�ҹ��b|W�W4=d�C���a9k�j>w����[�0ok4�n�d��I�X�m-���]����řX����q��X�Y!K13h!|	E�s��>��^�����[�s�-R4k��-���o�<����\��X������g�<�,	��9�tf�Z��y�͏�x.�~(��%$��������D�́�,oL������@j����^�2g:���缙�3Ө)~4�f��c6�9�k�,x��k�L�Ο/�O>��/�J�'�F�� L#��,�����31c�o	��m�l��d�.��s����O���/�����s�Fyƞ�L?�T���7a�+\���K��.�\}K#C�&Aa��5�6"vc,�%% �Z�zX��\~����(�-�ڑP=���*av4�a7�c	����q�K3m�J_O[3�8Z���
&�`�( jm;SB�	�̠C#X{�9t�FA�ct��B�w���a~QI�`� [ʆ�iI,DA. J���	�j���×NT4b� &��U�Q�� T$��e.�
�BH�P�i��Q<�×�@'��6/���x���Ǩ��Иmm��ȥn�X���N��$I6<�r�K\�2�A��Ⲓ$�p�L"�+m���҃�L`T�ӗu	��$t� �NWd6F�6�#��+��ƫ	��~���0?�p���q�L��>vHh*ƙ�o��wp���_�So��(,r��i0Y�SB�ђ��t
&��������8.���^7Kɂ�(}%"�6�(}=B�eQ�A�O�PE��Q�AD���<���Q ��;1N�
�F��B	�� Ш�-�)U\U\�K	�/gLק�vb	�R��/�}��>�J����>�~_loY��"�JPɄ+�f�$h�U��!
���Pp�@�D T���m�d��8݈��J�!��)�Yz�ZQ�Y�F�*%���C��L$�2�eM?,�S��=y�9P��m���G`�BL𲃹�LmL0�p�SW����!L-L�dYZ[`��9�!4�,'b��d��N�7�7���N))��<���/�O3f�P�%W�t:�[3�>� ���/O�Om�����Nvp�䄩|gyNsWJ�M�\&OT�7�XB��$ *�P#�
�ʰ|���Z�#�k�Ҕ����Ga��ɘ��s�|1u�D~��`[�6J��#�M�b�ؽ�\�,�Ր����
l������JB��tm����ڏ�˻Pw��x@7K���Ԕ�_����0,e�	�J�*IB$}@kQw�-������G�uU?P5�f�������!������>|��2�YpK/��O>$C���[ �T��(�RA�C��4Gyh3��f!�T.rO �t1�A�� t�NI!]����=8��<��Kx����}��y����ְ����1�FI �F/Ŋ���^��a��:�#� &6��P\��֝�8tv/�]<�{o�����������������G����7p����5���ݸ��e�{�*�+�)�/����B,&^�פ���_����ː�R�}O��_>���{?���/�{�z�����Qy�
�y��x-Jx�OR,�4Ȥ�Hd�#�!I{��h����n�B�=@���:%�$ �cO�x@����:���:��W�e�ean�r�I[�ٔ@��C�O�!����������l��avi�j,����`���v���=����2+�Ӟ��Ek���9�������6��s�*��|J�%Y%	Qi8VU�(}T�)�F4l�O�8�N�{�4d�E�a��w�ĕ�PԐ�hL� �����,\S��b@I2"%W��.�]��P��<#��50,U�Z��UјP��XВ��ˑx��{�� �'i]|��f`��=�/�|ımS[:65�`c#?�M۰�a��6bNC4|	G>������H��#�#!�qJ��Uu�hl�W��m��h������5�4K��Ų�uX�=s��`6�3�~-|�m�bV_�����>�����}<+���4�}����p�E���o���0�"�?�����Z��%Y���-fff�l���,ٖ��1%qbNfl��M�4M�rO�����WR�:�w���s����=3{�����z�{�(ɀf>�	+B�r1�c����S�����\�#�g��YD#c���2Yw46�M$q��!m%��Н��#�B2��k��E�4���e;��jo9�	@w̭[����yn���(1AT߶n���򲙹XBh���sb�D,ѹ|��$:�`1!�r����8,���F������L��7�{�4�]8���c��~ߍ�31{�I�N�GN�Cϑ�*��oC˞I��A��Y�؇�Ǳ��Y�z{����.a���8���Ǯ�ԣWq��8��y��,v�?��c�1�'���0���C|^�<�C��Á�����|�+8t�"�?�u�s�\���ob��g����|{/�®�'p��}8u�y��^��.sz�~���Ӈ�:3���n4���}�Z��e�����45��G�p'*������աh+�����YU�(�����F��P�X��Z��ʑ�g@Q�ܶ`K9��Qް�եȪ�@qK
�j�߸���}7�u��[���a�����Q�܀�֭�hoFA}�j�#{3�>kX�n�~8�[]��j�y�ʮf4�t�q�[��چX(�AGj��Q\U�"U#�0�y(�L@��!5'�^Np�����\�QS����[��L��CCw-�i.U=ݮ1ׄ���%@5Y�[Gp����j�ί�'J�9﬇�FX�#YP,0Q]h��AfXd�z�]j��ah����V��K��To����s]�`��	�sAD.O"�R\�$�%H����dЕ���\uW��k2�`T��B�T@/#G�`-���\M@���k	L��0�N^_A�.㱗��&8�D.�#m<�]���X�OTô2k3��4��3��"� h�bq)����%0����dC��ł�FN�𵵒��H��\1t� ������?�����A�D�bM��e�y����"\5�Q�d�WF!�5>���ๅ�& �99c��\�R�{��9��N�T\>C�h1�*P�zJGDŻ��r�h)��2��A;	X�xז����2�����P����v��߹I���h?�eHt�s�o%z��.����+Qm9Ӭ�~J5\T0*ñ�:��+8�z��z0��@��N��辗�8F�NAz�U=ݲ�/�l��;����Y�|Z{T֮�L�O5��L�jc�tA�=�h>OH�7��k�1xn)M)0����.�.�J�UX�~4�����#<���ZcC�Y����N.pt6���q鄀��/z#P��������@��� <2Qᜆ!4<^�^D�6�ѱQ���FTD(7�������'@��N�"Te*���8�u�tQ�O�S��
BePUw~(��:�А��T������X���
"t��r��]	]k=8�#2�ay��,FVW����4���6��>��7�w���� *c�6�?0�s��	@���0���q}�ʀ���B�<@7�lA�h�w5���4@���S�
�2�c��iL<2���� z��C�E��*�JO��]�7��G�@_ (?�\��3ئ �StǍ=�ys?��|���鎇	Ї �}_ލ�7���qR z��r}�Б6�
��Y�L��Upy��Eh��h'@�������H�4=܏��ZG�p�R����]������~i�}��u"B�!��<�?��o܇7~�6~���ο��ko�����S�����u4�C��3��I�����P�Hd�"��Rr��΂X�*�0���7ֆ��zN�cd�#Sc�֣�!յ��.�AD�/�R��\����x�G�9v#�=���k��TN����W��o?ě��|���\��s�q@��i��e��U�x��(��Z����#���dv��HHVs���@�Q���CzW�ܘC�lC�r����_� ��ձ;�)��#P%��z��9��;��Ghv'!���$�";�ܒDx�-)�lO�?�yg�&#�9>���m�AhG*��Օ��e�ٞt�rA��w"�x�ЁT���"v8�Dk����97���ރ�O�Ɩu(D��Pİ����HB<�DI[Ui*�p��JT�zP��=}�[#a���Dl���?�O�xO�p}�k����b/X5D@����ħdB״'buG��E:$Z՗�=�Л"0g+`�g3��C#BNs(Z��Qf2Yk>���!R-zRaՙ��86Eñ>6��0.�~��+�aQ5w���Ԇ�XԅaC�L�#�B�y���	�p)����hϙb8pߖMܦ7	D�'��3�ϩ\8�g�������2�o�w˂u_,aO,�l�W#��V����M0'�����"��;��@��W�c�.S���aL����ZW�
ay�G*a|������ kw�a�.�~��b��\t.�d񵃱����N��;C�S�H�]�#�� "�c�o���p�����\ˉ�5{ʰ�]�=K��%�������9��S�s��I'���d2+��W�Ph>ӹX�sn���W�]4���@
�'b�x:�pݚ�4���E,د��S���`&B�3��Z�-3�:��n^��מ�����~�1^��C<������������S8��#8��-5��Gq��pߋ���[/�ֻ���ﾂK/?�3O\��go�����=������g�����>x]m������?�G��
�}�	���<�������ޟ����s������}�?���K|��_��w_õ��3ａ�?y/}�]<��[x���w�����7����s��ɻ8v�~�ލ]N�����מ���=�˜���p��|��k8~�^��q�޺��W.`����~l;���=��O>�_ơ��`�=G���	����{�îS�p��9\�� fN�ı��������٣�:Axډ�=,��D��.�B!޷k;&�Ď��1u�F��衽;�C�wa��L=�mG��|`��.�ݎ��;1yd7&�bt�4����ۊ�n^U	
7�������\����(�En�k�R
�PRW�pX����D���l	Pg��c��Zz�Vo-֙ib��֘�@h�-=h9�C���5��N����ռ t�J��0�bP�3��\ h��i��F�Q�g4#F���g�����ce�3V	�e���bBt�D��t1�(�W��c=�i�%6uI�/	�6��+Sܱ(ܒ�t����$@%t�}aT���-�:7��2���tY"���/�dE�r��>�fU�j�~q(���}��.ź��*�
���Ot��9�ؐ��P����k	�U>����{L_>�/�;��7?��＊��ئ������X��ș�I+��9a� �r>S
��J���BjЖ4�Om¦�̈́`2�ʑ1I|r� Jt
@����*Q4P�L���,��!��wh�<@Q~�A-�y܇D� ����dh�9�ry�
������Z��T�y���˭L�}�����.�=U���h����!�3%���y�V(�v�H
�,{�G;˲j(�s��I�����c�n���=�'�����vq��G�ua��'�BH���A'�e����w��wN���'0|m
��P{r+�B�v��p	��[�q𩣨��C����L�h/���&��CS{t��ah�c#XX����VU���q���-\]m���Dt� 44 11�HMM@zz2���P�2&.	I	*��Pɔ��9�(������x{���ކ�k��Z����.�`8>]���/gxx;��ɚ�P}#]�W�J�S�k@�x�X/(��Z��XC���Z��k�a��r��^�Ekc���Z��7�	��a�(Dpq r�s1~e
�_��nm��憂l??w=���� ��ֳ]s ������@�N�a�ѭ�;܌ه��螇�a��v�� $��P'G�e��}n�݀��M�9H�!@�7�uBD����~�o��T�h�Y��cG����]S��&nm#@����G��y"��;��� ����;tuL�C.L7O|�?��K���4���c�
zuf��FpJ�y���`���F�]��m�c�����q '	�c/����q"g#��ϭI"o�7��1J�	>�"Rb�s!�f�-�h�LB�.�FM{	�>E��l���I�H�����B7U:�)ɦ��O�^"b���^t\�q$��B2��r׈.���~�?2�}/��_��~�������>{.A�@=6���.���Vp��G�#|����>X�3=��ㅤ</$�{!4��|�$��!{KR�g�� ���"���0�38�1�~�J�C ��D�:���%�aE)�m���q�ۏ��_�����
n�����^�z�$�z��ۅmO���1���s�j+P�vtK���#dh�N�>nis;7��mq?_Sm6�>$��2��E�Cx`��`���nN��7���!�)u>8���N5!m{�	�04���$��Q���HC��"�A"�cP���,�oM@HS��@�Kq>��!fCZ���<f{2ᛆ���s�*��M(#��נbJ�EH'���>��xT�W%6%�WȇW)��K�7��<�	f1v�4�	/��>��S���~��gi60�r�m���`̺2��%:m�В�L�ڎ�l���@�f�v{�y,��up�WG��%�iE��<��K`��a����B2Lf
`>��q�m"��^w6t��`(�D��$7S
K>H-���ݻ	��6����!
�l�ݱ-�?�.�j�~��'j�w�^7��`\.�9��<O����;��-Ah��0>X
�#�p8P�}Ep�S �}p8TG�Z�q�v�8%6��_�C�p�98����*8������M0=T	�����[]�	�S�`�Qmί&:W��"���mұN�?ym��ǒ�o�b�G�N��q�
�����3����%�0V���n����<�hVLec%_����,,��N��壄�X�	P_MG��j/,�&gs;BurȒ�����
�N	�~r�*{ڗ�U�}����I��oD�*��t�Ğ�w#�m��~��B�1'�eY�ib᳿M}��>��]S�?��G�b��8v�=8~�Y����;��O^:��gO`��ػC;&�;���ۆ^�{v������>�:�;���{���!�<G�q����}{��{v�s�<�b��c;�����)��N`x����P��15���hc�`��;'ѳ}#{�a��^�؉���3G0{��c�����p��)�����8p������8N>xG�%0O���>����0f��>��੣*vُ#���=�.���K8}�9�n;�����f1��483����5�ѝ���3v�mC����q������ցN2?8;��}����݄e�$�C��Î�1�����۱}�N��BcgzFY���¦���nBE]5J�Y�.�GNi2s�O�4-?>�~��4���#�	Ps��A��Vm]mhnЂ.��M�gf 3�1Z�u��q6�z7�s5�WC���jg�">%V8�aw�|Ͱ�_:!2�"�sѹ��TS�b��!Y��Xaq��̵]�u�HⓅ�1�*��9�X�XJ
%�T2���S�|򹿔�\��E2&h�tC`X���2��%���yo�cy@bm���R�WL��(LJ6s]���t�#�%z`Y�V���^<w,O�T�d~q���pˡ&��c��;˰:��,_H�R��J���E�XMd�ɟ�r�Q
͂��%V	G��`��h�s�n�:���^�o?��Žu0�kI���	Pö�$@W�3��j��^0��#垕�p+�oy4Bk��5#e(�Հ��Z>��:\��1�n���r�-�v��|��z>sk�7S��Y.ã�Y*=��L��gr�,a*����)��B�ϥ��D)����l�/�ϱ|°`�T�-�9�q�|�@��i޶*▯3d��$%�%[*���^���}�򙸰��#����$�x��9]���B�O�|V��<�u��wQ�g���6,��ߘPI�N����g�,+�����dȺX���#�@���o��igX���h=3�V³��\�]`�"�W��Y�&h���S��|�ͧ��F|��'6��$D:0yc'_>��c�d����Z���J�߰��[-�u�WYc}���܊t�6�R��>����D��/����@D��!519��HIFB\�rX��� <c���J�&#����rCxH �����X$�F����ħ���+�$H�|�UU[�����D�����`�h
3�����6�\��GO����ؤ2D�:Bt��T2�2f��*5���k����]S;}��!�4%��Cˋ=�b�1>�h���h����L42nO�t��|{��f�\Ȉ
>�*������az���F�NԟjG��64n�̵�8��9��j��F�~��;A��%<�;R��=��r���cu��p�I��z�m'��q���e���=q��d7��$��� _�[Q�����0v=��O��ɀ>6�ћS�п P��F�%��u;��W �v�O"t�Çq������|�]�� ���#��ÐaU��m���d9��N�\��e*�������� nh� �,<�S�n ]�P���:���]�/.���������䏟���_�����O|��_=��=ȫ͆o�'���t��yl<���S�9ܣ���w�1<#�a�oI�Z�+�EqMz&�1{l�����vl
uu��=�ӏ_�?~?�W�����|��&ξG^?�]��':������
�#7�1DX��w��?��5���P��g��ﱙ7��{�հ<�!��aW�h��bF�����_(ש�[��>X��GPS���H���\�5�3�}�Dgr	��=�x�nVUw����D�z0ʿ����= b��f�4�.b�Ѷ(�.�#/_�[�­g��[�gX�¾.
6�Y0nM�~s";Ra�s2Ȇ%b�<��@:��2a4Y ���0�(��l%�O���X����[`���;*`ˇ�ގ"�,�1�l�f�
`��m:���\���|�ʰ�E����s�y��;��S
��*aG:&	K{���X����u�9Ro�������C��?������D�S��*�����&�I0�3��1�krdL��9Ò�4'2�	X�Ce�:,ۖ�����|m�E�!8��-����'p59�vW�����\2�����x���K	�%�|����O���<Do�8��'�����my����k.�IFR�P2��r�p_b_��m�X:��K�Yn;��`*�����#<w���u������\hfbu/��I�rn�h��D�L��ic�D��}�X�c�U�E��Xf����i9B���,Do�oJ�3�P����ښb��z�5І��.�X�p����!tL��kn#sfְ��#�~�&�:Xk�����J_�YZ,�׳6���֛�C�TK�VcѪ%X�B�r��j����`e��_�^^_�E�aѲ�X��
�u4�B�g�W�R{�Z�4���5˿�^�3� -�ć�e�z<O}ch�N��3K�#�nlg�z��z���p���T�C��V[��:
b&�f�q���̌Բ���
�����&���Z�[��0a�5;��W�L�L���
G7��[�ci�<m������&�ٺ;���o�z<��q~��&#B�����#$:���HLOF_3��wec
��~�׭�g1�z;�l�aincCh��z�6hJg �F�0���~�L4�DwV[��f��4�Zwc�a�v3�jQ"�]K����y�Y`u�%��+�T���1��`�S�N�;)
��� |�Х�$gRw�T˝���4U�NX�`�E�2�V��B��� 6�I�tOhe���j�A����#"��ہ���X�ꁵi�� 4���<��󫓽���
�� ���^~(,+�aS��a�X�m���XK�je�C'/�����t<�H���vq��D�F�T��9�C#�k�mP2ڈ�\�C/?��/�¦�VF�1�X��s�h�V�3@5�<a©3��[� /�ӫ$�[�pe���(��H�� k�
��eȚ�rJ��I�3o��|M�E�5*��L-ٽe�PA��TeA�,0��F�ĝ�Sb�%�~�X��F��2H櫡\��N�n�O�rYP� Q�P.�3^���\	�O����@�9e>s�Y�ʑ6Y4P�ia*U���m����TnN��Sd���<�&C�<������,?��TM���׷���8z.����zΏ��� ڈMg�<@;���(�)�r���^�;��L���z�5����\��#�&F^��uԁ�����&<ת�nx/3�=���J�����LN=���f,�c���x�1ш��$&c������
TTU*|f�)����<\���̦�bd�& %>!~p�*�.�*�����;\�d�[�鐧�!j+[������04Ӄ���7W�Љc8x���Y���$�yo$@5��N�����<�sg5�]��Zz�a�n��� D˰C������<���=���|��׵���<���+ ��B�\���2�[/t��ԝlCݱVl=�I���ѧ�`Ǖ}8���Qb��;Ђ�m��3\����@�l@͑F�U2��
���<M���β\~~PeA[�w��t?&Oaۑ~��#�vuН�T��' ��@�O�~N=�]T����O��yo���@�<|;����vt�����'^���/��q1z�ȸ>�����۲� ]ȂJ�[5��B�%d,ȅ�9�.��#��ޓ�¾�
P�ޖ�Lh�U�Zz��1H0��S7g����8��)\}����;���5���?��{?{O��$�{�>�x ;���
��e$|�|�͇�}�=�|�`l������m�������ݏW?z_����?�o�ߏ��#��ś�����������C���Wq�{7q�s8��q�~~v<�C�s��q�=<��G��[26� ��d�{y=|U%�����>%��:|��W��9/Py���?\B5�NE���."�+Q�i��m8a&��W ��^�_xM�wF`c��ylF8#���%~c�Rߓ���4$�� m0�EȞ(�ô|���$`�hB�|hJTjDžZxU�8�fQ�(�,ģ�<�w>~�>{�����f�|x����#F��q[*,z�`H����3�J��y&SE��.����y<�C�!B}�0�>�D ֫�6|8Z��}�0�I�n/���Bz3y�e�*���r�
�KƳ&�J��Bs���JX$m���Z��c���@Lx�<G�X���v� CE��˃i[����4'�x0�,$�%d�\�=����϶��ۋa��<�־Rl8\�#�� Y�C�0 :��I��<��E�Bp^_�����dA��C�蔬��Y*�����i�0�wƷ�92F�bU}��z�
�Le��B���b�x��t.�T�_
:������r�&�S��[�r�h�����O����u����ĥ�uYW"��EbͦphTGB�9F�������� ��tyw�j�������P��kc���-7`��.4m��AIo���N��B ���#�G���'ԤW��U�cA9BaA
<�>�@�Yi���Bg7�G00:�����CAi!Ҳ�	7@X ���D@�Fxs>DQBj"J��P\^��!��%�Ӓ�ra�~s2�_��lNc���$�R�����͛�?��EO'ZZ�QXT�̬tvw���1�Q���BϡjS%�K����u���,��!�������q���DqE	��Q��SۧT�>Y�V�G��Er�����*ji���"�#�ʚ
ln�FRF"�cÐW��MuU(�,Bay
��[���/53�9��\� u�||�k9�(()Ė"!?[]O��r����AD��O>Spx�X -@ҿLLN@v^6R�S���r}R
�mi1r�s7wW�K��^pr�����<@e����76���6�A�`=V��"�%XA��I�'~V��6�Z/S�a��4Q]�f�fX�iMs��U-�<�K�P,w��3P2�A�|t��	����˒]��Tŕ6��ӥ�[W��t91���5��aP��"Dץ�+����c����B+�@��Uӵ�O�ZGdjgm�nn04ӹA)�:���� �n]�7ք9c�??w���C`�����d
��}�s]V �p�k3	��`�oĊT_�H�tR��U�n�Z�L�����~O��"���(���.
�R�V ��x^E|j�z�"' N%�𬌁wy�*X0ߒ��&���*P�g+r�mA�$qFxJ8��I�M�p,릪TT Z �q	@�T�pJ�D�R	�^ɂ�x۹����J6T���|fL�@�ڤ��!ZJ��T��� ��TA����-�E\*Ė)lގO	Y�zЕr�N~�Y�h%2�x|>UF����t>�����]�=ӊ�Ƕ�1�n�X�s�ؤ��6���X�R#��$�>
h�o���9�>0���'���;/Up�>b���8;�V�
ɺ��G��!�Жs=,�u��|7C�����C�p��4Q� s�6]��X���|J��w��cv�>������pDr������d��7�������!3=)�gfz���_��EE�'7oތ��t��>������f� .2�Qa�v#,	P_O7�;�N��޼��I�CD�����u���v�氰1����s3�m�,?��)�o�Atb]\�od�uZZ�:�z]>�4�b�dA��Zs9Vk-��S����E�U���R~�����x�i��\�yiH!T *!�w(�3� T�a��wW{��·���'0}�N��C��~4�D=Z5[���R��7� ʲi�ѭ�?�<����o�����4��o�X;�N��|���EmA��>�[uB$Upg��K���6t� �j���� �& ����E�W3���v�U�2��������s�0y}
���� <�g?��O����v���M2����˹(�$Z�����j*CyH��op�?̀ʴ�[Ur��]\G�m�[�'����wc�{p��c�������[�x��׏�����?s�O���?�-���'���Gq��p���{�I��������8��T��{�#�/�����x��G�T���*.�q��?�}2�Γ;1��Nb���c2��$F$���(F����>�<������������[ |�T��d���C�E����#��^Ќm,��Ў$����h*mA��h#���>�����B�nNP����D��Pd[��>���ԓ���t$d"}8E�_��-(�C'��>d�vU��(��W�l"խ�F�ְOvŖ�ͪ
�G�=��^<� �l��H;R�H�9��y�N�%��U�p�4�`][<�v$B�7F��*�i.Un�p�&P%�i��̨dA���8�j��&���<�KVmGw�@oG!6���Ka���{�`�m�T�D(��P5L�VL;>��g��<I�b��(hn����xX�$á.�i�j-@�h-�'U�0�����չ�/��p��saҟ�°7��x	�xM�w��᫽����_��,�ѩ��x�W���~'cW>�AO��G��K��۝�e3RM��&�&	���Z7%�3N�(ayg,� ʾ�^�(�-	�1�@r������"�e�ߪ���E]1
��z��D,%$0;���=���ZO<�KT�R��W��E�¨ reQ����)y`��1�YaI���UGW����x,!@e���������,�����c��V�0�ԃ��6؛A������C���F,���Y�#�DVAWD��dEe����}�p��a�ܻSۦ0�cG����W��3O�g�������˟�}�{ϝ���)t�����ׯ\���	~�՗���?ů�s��׿�~�|����̓O��g�Ə>���o���~�k���/�_�
���Wx����[�����x��g��C��~��s������w��>�_~�{��?����k�6�޾���T����wq��u<t�*^}�%|�՗�C�׿��{�q�?�_�xo���������
?��'�����*��أ��＂w�}��]|�����~�������o������_U��?��O�λo�'_~�_�������˯~����߾9�G�����_��Gx�������K����x���!_��'?Ɵ��G<�ģ�o��}��ŧ?��?��5ը�݂ƭ�z��"0<<���~S�۽�^����s[9ާ�~��/���ط�]M������,��^�J�t�c��6����XnL��.�
km��YCo�-����o-?Kh�2|,��m}73�s��
�XᢏU>fXH�[a�T�%2���b��JUܥ��o����qt!�wP�
FS\Oo5��1� Kw'ʈM�S'�Ou<����{j����K����i^*��9:Ҧ� &ő��J�]uLK�`�e�M�p�I���d��Yi4�I��(�%��<�����鬀��t$M�¯���|ϖ4�N��n�.u#?�'V%�`C^�"fZa�Fk��wP���嘇^{
U���u�n�'�3���}���o9�w���� ����0>���s �6	Q��ș�B�ޭ�`5R����s1�U0%P�%����v�O	���4Z�m� ��U���\���@Q�((,fM#}�@� ����M��x�R�v!*!C��oc���v�7U{eH��,�ݫ��|���s�й����i|VKF4��<�������c�䓻@�̀J\g���Җ�=�����Tt��_�����M���It
<���.�S�%*��o���P+,w�9m,��ߜ��G�vG#�%�n�
�W`��
�k)�ue\O-�������Ğ'�����
	ADT$�	���4�3���@~n.�JKQ^Z�bB3��Y����&@�A�����Ũ��S8��X|�?	���pr���=}����?o��)�JP_�IWB�v����]�ajiO?t�`ϡ��iڊ̂B�VoA��<�l"��F��"@u�Cs���b����R��X�~V�_msM��9!���%������T����@�e�����J� �z`X�]ȄJ,�]@��w��}�h��a�|X�v��g�G���C�4lÖ=�(��@�t�h��&�o�����h���Bt2���C�m �>3���=,�<$��Na���}���H�O���]*:��z]�>��~��{	Ѓ����� �,��{��A�x�=K�^#@�2Jdܐ�W���l�T�2����\�20�����C�Hz�y�W���I"t��#>�s���������;�	B�����˲ T�����r�_Ug&�F�c��m8��a���E�|�&���Y���7��o?�'�?��W����	~�ߟ�'�)~������!���O���?�������C|���gd��>�b|��?�S?xg_<�3/�������s�����}b�L���M��y�P�Jȹ�T��J{پ+�f�0�����_zyTt�
ϟ�#C�\�-o��_u:�}�G>�L4�7YuB.UpۓOh*H���"�%�_h����5aM�/+�!|��!(i�zhS<B[���DD�Q�q�h�Adsb��Е���T$��#u �h�h>r'��;^����ܳy|踕��"�K�г���)|���x��>Ԁ�|w8z����dUצ'���ɂaW�4FcmK��`<���bXN��d��-R���^���s�rQg�؞e�=�}U�'$-w��%Z��0�U��U0�Q{*�3��&X���l9�����#ky�47�@sl�f�����1�����x�7���^��g!����_}��~�5>��O������	���aZ�,�����2�U�0��ǆ�xhU�amU,̇�`��g���x��	qlt���,%B�{�X!T� xj�)$T9%R>w�a�4AHL*p2-�+�W\��-Or[���X2��� *e�	i�9WM��!"e��P��"1?��!�S�)�$$eh���'?�����^�N�.�&Pe��i��܆�\җ��=�XQ��lTgq�K(�j��{hm��FW
���<��"鄨��'D�Gra���	b��d-6�n���|�YCO��hE��B׊�������)Y�����+�DF�#11^ecb����v��������,`onw{$FF"+)p��E��Zj�p��9\��^�<xO������ѽ�032���6��7�iK6��(3,��䢲���غy�kjй�	��ն���**Frt4��CP�����Mܮ��IH��Fmy���1�Ս��6u.�՛Q_]�
��

P��Ug'�������eeH��EVJ
���Q�����r��lF�j5_V����Ҭ���c#C��,EYI!�6Ԣ���=�n3j�lBC}6WW�m��H9NI^j*+��Ѐ�<֖�
L��N�MMhf������������Ņ\ފ��&����G{;x�������6���Bey6o�BZ
��a����P�f�&չn��������_���{��Ӆ��P�^����5���QU��,خ0]��ƫ��n��~��C��!�����%Hu�m`�km[=,5\�E:���h%�8l�Z?�	�Ɗk,�V�JU[���"�K�nE��E��ХQ\���ع6�!]h*�L��r+-Oq'J��"W���j�L;g�j��:��14��a^06��ħ�a����d�2�zĩA�FF #f��,��iQ8l*��X�w�s%<���k)�[E:�r�a��M�p�LGT_*�� ���=�H���-�0ˋ�Cy*�`Q��0�M �#����˽�1xf7>��_���|�{�����J��:1n<O?5��
i�JP�$>�%��:?�D���_����t��%#� ͝܄�M
��#%�d?����BPY'�I��lO���!�)�m2��Nɂ�I?���6��(0�NB�s��SEH��d����@S���Ȱ,�e@B�,�Ѳ�uj?Ҏt��л��|.TÝ�<U������2���#,�?�C��g�F�5Ý��:�y�d@'���5ɀNa�~��	О����g����$�T�!t�R������`��t��7w��� B�{�s��
�%��\���+�Aw�7c{�������t��� �{mL\#��q�OL�<�T��S��`)Z�{aFF�z-5U�{�"�����d���ۥ$���	 l�����_W'��6�ư33��	���v�����+��w�@?��^�<G'������ ����	ޏ�\��������PR\���T��&Ʀ��� mm-~vMhi�D���j���떫��˵���A�ɾ���AXy"k����X����L.d2:����� Tb!*m>o_���.�nm@�O�c���q@����)tD��V��kA����p�5�P{���k!@y�?݁�3�**�q�G�m=�8=Ww�L?f��ˀ���8��4f����|j7v���s��m\?�جʂ�KGD����줪%:-C�\�Nx��ץWۿ�s�������1~��<~�=�}Ş�G�SNo��7ĉ�Nc���o�7�TЁ��BoςJP�6�F��J��>��?�����(l�-N�E�y{,d@o�~J���P�3�J�
B�$C�h'F���]'����9�ᛃ����2�Q�f�O`�c�p�	wg/>����kuG�8D���7����}oߏ3/݃�Ϟ��gN��sg���_����{x�'���_��7�6n��:����7���a�q:|��#��e�(5��|H�X�Eӧ��{�[�/C�܁O	���!��θ6��)�Ioi�r��Z�N˵�u��niw��ϱSs�"c$���4���X *7��[U�|�1�w$�p%�ޖH���g� �!�\�J��P�J,�S��J(x�
�wh0�)�k��[�����#[X0����HF��ضxB4)}�*�{xS��P�E���FTE ��K�7,	P4����[���#OF!�b�7�W�ô.��D�јX6iO�Iw�@�|}G�xm�G�T�C6���t4Đ·� �0/��`6LF������p��Z��ۈϙB����M��ςNo&��s��S:#*��M�Щ��Ss.�;J�^��>h':�x`��V��/���������������_�����.�}�Xx��>�_x����w_��g��`��Zsa]K�n��eo축5�]���!>5��AkO>t��{��f&K�S�j[&�H/�۳�B�h���;��s�h"��	����6t.#G��F��n7�b,Tw�=E��$$��*4
�q� �3��Œ�����e���j�;����M�ډ,H�r�t���쌝{MB�;c���}m�j�ε�QH�Ն�??��7�_����5���,ǆ�T��>	�%�i�Gw&�j�&</O#�����z0�0��jk}�9xJu[C�����X��BT&KO�Q�,4x���v�V*,Y�06Ї���hC_w�t�:Cq^s�*�X�kW���p��m�and���j���r�,_��Z�050Pa����빏�X�b9V-]���ey���6�f��ֆ��>ܝ��dk���x|{{�~��%<��^v����FLx8����|a��#�L�his�����Njy=��z��Y�T���U+��vt������o�1̌��hg����/�~&�\r���^�u+WBGc��F���ym%Cs�J�kiA{�hq;3=}�y;ss5oah'^o��x�&��uՖc,_
��������;l�,ajls�K�N~gF�zX�nV�+ym�x������G#C��	>ޞ��򀕵%�7�Wm@5t4@u����t��d���4��!N0	s�y��a@|�l$J]Ma�d�Дpdm΃OR�Z���k$`��VXf���2�t�9��ay�%V�۩����3�QɈ
HWF;@#ѕ(s�&q�>�k��T���UI.��������@�J���87,�%Bz�a0.�"4��3�`���(�´0zħ.����1a��U�u2�'Be�AN ����/��A0"beٮ*��L�k]<�2�P� ��txVgS�8W�D�f�1�n��3v?��է���d��#u�	�up�N�sY",Ӊ�HO��ƛ�����s�|�q�����P�$O�!��߫	�U��h�NE��MEDC������;j�5�I���h��h51X�B��\���+S"T�s.沠�D)�M�e
���tJ�s���yA�D!(�4d��������kU�DՇ�Q�_��4���VT�C��G�Y��Ǜ?���è��K��٬�ڦ�Y<��p�����)�H�C�H�v��T3F݆�g��� T��h�8��j�T�+I��A�f��ݪ������2�2��vb��:ϱL=�����$q$�#�k�Q)k3$Zw���%F�ޅ�{'�ܘ�@k��hc�!�G�kx_Xǿ�
�f��;����쏰�P����iHLNB���H̥`s���ԡ���-7�-AU�&dg� **ᑨ�o���*+*T�4��%��~>��":���� [ؚ���.6Vp������.N�	D����(��!""^�Dk�;l-��ᄺ�z=}7{?�f��VTl�CCc3�;�QRZA�����|&l�3H���u���~֬[����b��eX��K5������e)�<��ɨ=Ѐ�Gfi�A4�����ݜg���˻�3�;C:�A��l"@��T�����>RW��2�u�g��r��bە=&@G�Πi��C���ۊ�NT��oU{�QwD�^����B%� P�PF���>���$@0}fc�:�Pɀ��,*�)uķ}��d@�)�����v��6���qM��܇����'Da�#�	��8F�&@�?|{o���
��	-�:σ�3us|����^p�*�����4�u��+���B�R5����'q%���t�sэ��s��������#F�0D�r���^�p~��L��4�3���bǭ1�>2���g���Y�yz7�2�<��ޏ�/Ǳ���Ӈp��8��Ic�{�����)�	b��!�W�����ː�N����P�]�� �*���k/�O�ǀ�w�N+�~�.��&�/�n�� ����t� �BF�͜���������#B��q��P"4\��2�Z$����y4b������x$���)H��Mx>��S�=����|T�V���b8d�+�֍n������������v���p*����UGA�*6E��06�̀u.̈0��Th�|V�<�xl��b�J�p�8�,�q`����#0�2a2����l�x}mw�aA�Z쬀�VS0�/����ܿ9�n��X�6���.��Y����㻿����gx�g���_|���'������/�ӯ?�W_|_��|����{o���_�K�y
/����Ƴx��W���/�?|I���������O��M����͗���BX}.|�3a�9������}���۠����K��� :;�=���S�7����X1���S�9IDJf�_�8:&Nn'�!	OP����LĒ~B�[�}�����L2���K	�%�	Xҗ�Œ��j����l淂�w�`�d<�MYn���^�[7��ń�F{,�I �$��d�m��lL_;�7��|�>��?���x�߁Oz8tR|`�5	k�y~|T,�����/�y�X$��X&���!�mL`�0�%⬉Ok3Y��001���\X`pwuQ4s&l--�@�x�K�b��
&Ě!��)#��>�)&0]����f&����A���Z��\�^@�s����1,�MU�����pqr������:{;8�۩�p�zWWg�N��md{��Ն��%��=�ҹ��B��m�c8p�8���ikk�'V=�Zg~^[p�Բ%��5�+��"�,aYv��ޅۺq[����c�Ǚ@����=�mcf[S��x�uua���O@��:*hZ[���s]=�׆1!o�k,�ӂ�d�g�y���t�^l���5Y���Y�,	l�-�^����jٚ�����x_�f5����$���A���z:��oC:\�1��*c,�[�����(O8���*�F~�0��������QӺO�����Wx����8�mc�t f}-���D���<�+7Zb�+�U�VXb�AVXj���XI�F;b}�+��\���kc����k�T5Mr�F���:kT�BjQ�rB�����J��J"mQ�-6����MT�M��~��`D|��%��!�[M�r�T�H�.��|0��s;���eI$lʢa[�ª4
��qh:�x��Z@|��<7�١p#*�J�a�	��08o�3i['�/@�A>O��l,Clw�������}
M%h���[?�.>��<��3(멃A�t�ym�����0�~�&Û w�:��H'Dne������>�R�Й�:!ʞ�çdA%�)�^p� *����s���pKYH�:ب�K��~J��
"u�
����@�j�ұ�7 %�n�B����˽��S!���L�L%*�쨠�Hڟ��Ce��g>*�l��o>*mK�P��v��!A�L��%:Pɀ�M�+�֞nU�ϱ�w��<�zĕ����Bt���y��,SMܚU��6ò� t����j�2��*lJ�A����m�{���S	�l���ԟ����^���[��;m��_	-�U�ݰ�4ajH|Z��|<��D��c������tO��74bﾃصk/�[�	�<��g!''�y�HNIGxD���PVV���N�!C��&� 9�� ?z{"��~R�V2����^k�{�/�!.���~+������&��c���hXD <��anm�s����/��>ōG�̮=�o�@Q�fԷt�҃�q��@cs"�c`"�/>���^�E���Z������I��X�v1�,��1�q�����DTM�G����<L{u�;t
@;XV[�Y��!�h�W�����<��L��!*��*��#nץa���A��nL�2T��٩9���&>��p�eӒ-Aٶ-�����M�?֦��h>�9��\����U�p�w��d/�Nc�@��*S��+��:���Q�H �v��z1��������vu����K�Z"�� ��qy�N<u�?��Ǿy��u��u�_8ł���|fO�e�����*���*��x��z�ȿ���Q�+�e��T��.�B���nN	Q�F;��EוnF?O7�׉�˝�ډ�k]��I4vaT�f����*�W{1|} �D��#S� �'n�aBz1��!�	�>^�>^�Dh��~�x#>�9�s���*?�^+��P�ǧ,w
>��Σ��k�ʵ^�b����B�F�k �?4�W~_2���H1b�T�%��4r��
@�	�6B����X��GdSb�X"4�%�qH�L$>��}*љޛ���td�g���WQ�U�`6���H����v�>rϽxW�Ϣs$��vp��metJ��S
�jDcKԬ3m�X�sY�H|�%�p Cyp�*��$A�y	��lNs�z��Mp߹|�:���o/"@K`��H�[��p�Y��R�T�C�8,�$�4!w�C��ϾK����?��d���{������~�:�z�q���Sx���;O���?x���|������w����|�~��/H�c���/�����K�᯿�׿�O��,.޺��ܯ	��~�2f��8�f�ɰ΅fW<�f�a����Ak&k&ұ�X\>���c)X>>Kǈ>�r	�_���ؔ|
8B��R%���K�V,��<��XUa��^.%,��+���.��2�L�t�b����6��D䷂�侖qߋ�ù]4���ܺ���P\�I�w�bY7��5���#�JB�6�'o\��}�.��;/������x�$t���!�kˁ^;�%�kzұ��?�d�֧�����XcBH诇��!L	OA��9m�UO��6��5���!C���`FZ��GJ��>>p%
�OԀx\��� A�'�FF��������D�A*��(�#��p��h/fp����K�^)���?�>�>���C�j��m�\ոvN2���tn�O���m���3G���֞%��3ʿ����Xx��d�p�����2�Li�ƍ���PYTu��D�d<%�������������)� //�Og8Z����uwt�+�iga	'Bߙv$VmX��&Reya�dx�2�+�4��s8����|�le�=k�NA�8�sp��0�B��w�̩�a+H�q�|%*�r�'�5�Y�%>�"ɀ
@7��tH%ðh���:SM�� �8�	�p
����-L<,a�D��[!(6���מ�G?|O��$:F;a�瀵V:P÷��@g����c��9��[`M��
�!��k3�:���y~��Ќt�*�/��j.�\6E�p`��<?���	�h!뫒�)6%q0#��2�������.���҃`��i Q��?���yُ1!j���yA�	MGއ�R�Oh&�)�k�D���D/6���mʆW}���W�ء-�*Ch'�;;�Qsz����m�EDg9�Ja�����G�X=A'c �!�!����w>|o~�6}�i���v��g�N��f�?V��ӽ�R2ŉ�/�oM�ˢ�@L{�	m�H�+B֘��Y�%����!�2,� T�s~i��H36ڪ�b��?%*��,�T�|.��n ���ʼd+�L����Ms�pey�㡹v�b�sf��T*C�(�· t�J�TÝk��������\��oQ���lPi~�wc\�ba�|�&�(/!|JRV{X�v��r#��W�0��\�������7��.���L�$yT�DX.$�TF��QGF��F`�#fK
=��a��tWBWW�:0��!@�x�CP�?R��[����F��tL:��TR��QZ^���^��6r}	���QPT���\d�ťD|A1r��������DVj:R����������H��FG`sQ��|amh�G1+���#�qwELD(B�OɆJ&4$���?ۡ��/���~�O���e��aԵt����աq4�v����;4���f�l���	�o���}}��&ѹV�æƚ5�$D%�F{̜������U��g��`��S4�8��A�bHM���� ]�r�t!#����~�_��,37�߃�s�znn�Э�8=օ��b�}
�c綡�@��v(����!o�;�P���{��p�ٍ���ǉ��h;C�r���:���O�Ĥ��@��[������3��U��J�
��(�z�A��9�J5\�k{���T z�8��=8��Y�x��:��7�)��u��I�>wSW�O���)�Y�;���>�@T�^�~�� �'d����B������������D/͵!UU�%[+h����%D�m����,]�!4{�u��1p�qC2���������)�7�����^���_Ɛ�\����%���[O�#�Λ�5��m�1;x=�u{�MK������>����e��,t������L��v2�����������o�VB�!�	��4�.��Э���qc������kM@|[b�	P"4�+	�=)*2�Ґ՟�ܡ,��0rQ4Q������l
�u����ѳ�/�q�|����EL_6��CUl�aVӺxشg�}���p-�qw�y.���/���l�� >D�K�|X��i���;�}yJMm��n��-��f�6|p:暴uo!<z�`�;��c;1p��<v�~����{�ޗ��~�������o��_��#|��7�㟾������o�ƻ��~�>��q���������/_�{_<����9��E|��+�я^��?}~����x���x�5�p�Q���Cx��'�.������%x�������^}>%�p(��iY4�����χ�L.t�s�9��uciXC8�%��2� H���
@>G������b~^ᓨ�'{�K����\"h�%��XF`.���(N��M$r�#
��mDeK(q6��;�m��	��ܯ�hV�cIV���YXCl�lO��6"���-�0ؚ��H&�����_}��7�}gN�?�_�KClp3�CY֗�bqyW�`Yi�KpCF ���@���ħ���LS��F�0r����5Ldc=5ޣ2��D���B�3%U35Ύ051�m�D��J���·�S�,K�q~^����ܯ5%���=aKh��`"�L�:�q\�Bm*[+��`�@#D�+;RU؅�t:�=�PA���zxͅl+8��<�=����]�Oz�t��$�����I�֍���oO�{V�*+,�s"�d[ik����m��k�΁ �̱jmnA���˕�v��1���n��D�/��{�T�(������r*�Fp�F��z#��W�ܕ��#h��<ߤ�D5 ��3VŌߗdM%#*Ut��%�*�Kڋzp��Y�tu������������Ă�K���}�0�1Dxr8���J���>����W��8[ %3���p��A�8}GN���X\}��Xs	������ߡ�-�{�C��B�:��T��jl��V�4Cl�V��-�0$���:�u��937�kS66f������ ���"7vż\�^��C��a<��Kx�w�Cǅ�'
��
��&��q�(�QV 6�xAO�At:KuZ�Ҟ��)��cE,<kS	���n[���Ɨ��(D�$�v���lAHWbF�Qrt 5禱��*���:1�r�>TA@K.ߟ��U����8�}�.}�F9���Dأj�o�����w��;/�ڳ#�����
w�v�7����R2���j�S�$w8�E�gK"\K#`�g�gq8b[���S���J"��@���܅6���R�|o�j�)�p�3�9|J�D�!�T՝됨`a(�TڇJлT�sUo	�y��E|nJ�[����x
@%�)S��W�'�̜���>l%*Um@�@%*UoSǥ��\��|���|�D��L�^p{�������˩��Te�H��Zb��$m�o���C�
���}��g�[ځ^�TUl�ͅ���g�==j*P�o�[�p����҉x��A�f=4��A�@�ħ��L�x/�D@�SbQP����|2�yY(*)b�����Am}��Q^Y���LЪM5ܦ�iY��܌��������C^V6�2�������(��s�x��uv@4��y�	������--�fc���z�=�!��B��B���`�9$<M�ضkM���RCtaxj�,k�mC;��lmEMsZ�y��Њ�Z�a=�QZ|��TCjx�#@�9ú�D�j��\��p	qDlY4b�cR���|aC�n���|��f��A��r�j~�!(U���+�:U/�����64� @w���#�L\؁�#Ch:܋�}���ހ��-(�^������Z��V�Mh*c������
����޹N��!@�C����x�?2*|��nN������]<i���^bt�J�
@>~ǟ>���]��'���GN*��~9�Ko]űgO`�?�m�G�1��4��P�mA��
� ����t�㜻��坱�����u��/ �C�s���5�^����y3h��G�|L;��n������*qE|v�=7�����Z���!J�M�G�"���	�k��^c�>����7�k<�U��J;���s�;�����Z�s�9��\�;��������p2�=�@��ߣ·ǖh�}�
��h,Q� �hAh��@#���V4Kp��B4፱�{턶$$�� ����QH�H@zw2Һ�����IE�@&�s�;��"�7yDijg2�Ca�ȂY�#�'���;�󟼄>��}';���\w8l
�kG6Z�aے��x����k_>4K��&4G�c3�w��y�A�2V�(��T�Zz����>Y_>(���t�C�{�x����|�������.~෌?�|����}�:�x�
�|�<��%�|��]ߎ��?}m
'����}�8~�(��®Cm8r~�.c�L��M�h��̶�|�h�����y����=,(�g�x�A|��w��O�����������%~��_���K���k8u����E�������0�	��D{�5�I�OǺ�T�&W�+�ƕ#���Ɖ��4,�W ��.�~8	��S��sF_<����X�F,Jf�U�ȐeTй�����s'�:$�1�΅hQ���-ܞ!�ՙ̃���m��<,���J�sm{4{򰴙����W����{j ��xꥧ�/qߥsx����W?��O?Kc�1т5�ې�UE�p�/E�Fd��S!1m��t��A[�� �1*�N��	��ζj�KS��X[Wf�
7�]�$����L���r_MA��T�I[P}���Ȑ�"=��*�H�k�m�y�z
��?[Bˉ�Z ��a��@<��TuZ7�Ο��6���������>�, �x�򺛧׹(�Z��V��T���R�d))5	��1����N2����k>,(I���%YA�-�f��!�Yy���6��%�.�8v�;������j{m���qq���;����Ǐ@���ӎp�jŲo)�q�aa!		R=IHo�~�
����6v�j�"���VY_^K�$�L(?�5�6���e�3���[�%߭��-,̰��ɀj��5����̬-`(�k�wd �@w����Ɲ��� Wgx���Նߋ��Cc�x��e��x��Ʈ]S������E0s2����}�``m?+h +@Կ�k=M����͠`�`;hB7ZcA�L�r�f�(�{�*}#lr�a���$O���v�a���Cq���	���}`{�?��}𯎃A�U	�Mq�%0ͤJm�?�s�`]��X��Nqp!6=x?��-E�`b��7X�Ȟ�� �O:�i@��&$�a=�l#���B��aD�T qrr��!��m�j������1εIp��1�+�������מ�������|�g_�����2hyYB'����52|�R��!@����ci8ܫb�Q�	�,R����A����YO��~P�����s�q�I�S *���5ᩲ��ec*�ף���`+C��̵�?d@e���v���.�S��NK��
��@�*��4�?m<_�K�+��y�P(�)mA�v�<g��؟s=ߖη��WSA�B�ܹq@K@+�ԩ*��O̢��d%����T�ey��a����me�}��m�1���,g��T0*�m%�)U�wn�泽j(Y'��{����6�^�DDu�|̰�p�lXm�u��j�PO��kDE�!-3	9�(,�E^a2�憅*�,GyU%J�JQ��
3;v����ą�@eu�Z��JD�%��o#:{�q��G����عk/{����
����Ɉ		Ed�F� �w�y/q����P���p%>�x�0��a�)�ԛ��@?o��'���y�~��X.DWo7���]�뽹m��؆����8p���8������.t�{l�5�a�{�*ޫ��BK_:롵f���5�`��
��53s3F`�F�m�GpEbZ�Pu�	�O�F��)�q�����oT�[A�7mA�1*SY�fYZ�s ��Sz��=A8K�B,wM]�I�T ��8��c#�z��G�Q>S�̾�����`+�wb�Iɠv��h;Ax�G+���?Ҋn' 8���^p�n�(d�>�K��OχdBe��W�U���CJ�����m�����o2��%zu?�y����r���c����Gq��a�u��� �?�צ������6�=:�BT��>4��y24K� T��h��d��:���τJFT�����%�ĖLպ�r��K�d�<,e���F�
�1�F�?�s����qZy*y���s�~m�Le$�I���T���n�L���� �?��C�Kt)��59&���G�ln?�?ތ��������<��.�=<�L0y��om7UU_y����v��?5��ڿ�W���@���$�ֻ�dF�����1�� �lW(U�S9���X���xc��N!>e�d�v�"�=��|`6��I
�ADf��xl$8�O��4��c C*m=#�}TCbycۚ����oJA�	Dm�ې���8��1g�K��6���X$5�#����"_��X$��r1Hl�ArKR��J�&�%"���nOBRw*�:��)��,�EY���'��?}��yv��,��0Y���)�ۚF�f��m˄U[:�z��ؚ��Ep 2F�p.��h9���%��#Ű�΂I[��%d3|w��y�.,̰���	��cǓ��Y|������~��_�w?�����~�#���>���?��Wwc��,��Br}8���P5����\��e��'��	h�5liKA+��Vބ�QZ��,g�������T�^���Dt§Ϗ���\�w�{��,���cx�+x��s�O�����kH�Fa|��9;��-�0�����qN"�G3�n$+�	�d,M�
Sb�X��KG��8�+&���!ç,��D�>�f��\<$�c1���/KeH�r��'�b��7v.�2�\ǐyU5��ؔ�y����\��ik8!ʂs�MD�d=%���R�M������+�R�1�	��L��;�hK�*��W��@�&�-�c�2�׵�����C���>�!��o�>�"�>�~��]|��q��>hj�a���=�0^��x��>�C��/�P�>~�Mc�X��ku������[�0�0���L�T�[K���|c}��l�A"�f�IuW"���J�5�v�:���%jutM=���R5T�y�9&&�scC�T_�m(Q3QC}XJf��		BPP |}����G��(|z��`Y�qvqV�VzI5W"U�%����T������;_s�L���>��^�Ɨ����E0���臨��ڍ��r|��d�������ԇ ��~-U��n�s{;8��zj���|���Dt�zy#4(��*�������r�P�e;A��ř�%%�2���v��<?�x:�s�c:�Xr>2/�]y.�%�M����>}����lma�B�������=�~�5����}y��c�Jkh�SCH5\s������cd�c3}8��#*.�~����%��w�;=�e�'N��o~����sx�g�ŏ����b��:���3��+��8����0񱄶�4���%S7Chyc=�:��	`Za����l�dM�Zb]0qJ��r]����`���K7���ND����3�z����<`� �l_Xgy�:��Y~0��)��90���i1Z�0ؖG��2
���g�7���1����S�~|&�6g���\��$v�acO.f6#��P׭I�i�6Yp�sͦ:�uq�lK�g{����/�f���zB��:�͑q �g�x�çI�_�ŷ^��'�����,�>��ɞX�ꉕ�|�2�d��.�ݜ _�;�-��糵3Y��y
w�x[�7Q���`�
�SUȝ�@��tH��;6�xw-�X�|P��̙�6�R� �W�rB+�nƦ����[�2�B+Y��,�@Te*籘>E�22g}�($@��ԣ\�Kh����HA�T��&C�HE��@*�:�� ���T�
@y��+YP���Di)�M���O܇
b����� �����V5��S��M�����&e��Chf���l;����h�s]�6��^���e"��(�.�c��iU��(���W2�,K^ bγ�vQ����i�i�O�a�Ai��G���Y��*��X��
�����G&��l�V���/�梢���hmoG��&�7nŖ�:��s���޾݄R['
�K��UjF&�x����7�y�}<t=�h�ڀM�yR"�CC���L�y������������/���n����������|y_
!^CC�������Ƨ�p��+h��%@KQ��1W�vd
;���#'q��p��U���e��M==�A��8R��oex-�K:Q�����+|j-�3-��� �*q���c�2k����v�]�?.�;�,�7���D%�����_��)��H'Fj�������o�6mt� ��l6�hF��F4�ۮ�®�����߁��c��ێ�����ވ��"MVcӞ��9Ԋ�c�;���D'Z�P�l��D�َ&�o<ކ:�Oe��H���a|'�?<�
�3�������;U6tF ʘ"B�	�Q������L��T��5��	Й+|��*���y� v�8�����C�q�+x��q��8q�8��8����[q��K8��qL�܆m���v�����Ó��B�a���,���L��b�}���P�K �?�n.@�ߊ�m�P�d�d8�.�%翕�c8y��7 e��Z���D���w���nqg�Uba��Cp� ��CQ��;B��������o��Anl�Cp!��WF�}I���͡q������(�*��>��'waۓ�UU]������\�����p�&�ߕ�hb.���L$�dsi�!��H>X7�΀�.�uQ�%�[@,Jf4�>���$��)�b!�ؚ��&�����������ራ�@̖p�2���d)�Ӥ�sK$�6G �Ӕ�(�7���ڹ���J�qDX1��PN}�B���Ʋ t�o��o_��~�4^x�&v� 8�	N)vpg��fK̫�`U�{6ڲa՜kBԡ'�����΅MOl����G����p,��X<&��ɇ�׶j�qމ85j/��( �`����-���S$ş�G�Ie���C|�ֳx�٫x�0��+���;7p����C;���Km"��x��ߑ�:b���OOGFXș�5�!�w6$cO}vC۫"1U��� �������	�ȖPt��1Ԓ�Ѯt��dbf��v�c��f>3��^?�����~������7��O��1�����=��m�OA7��bl��2:C�К��
�r;��)X2��E#�X6�����PV�dc�h6���%���P�d`u�p�h(y.�I`.陏�x���X���=Q|-��	Di�)��i��S����&ATr?㙈}d
���`�V�6��	Ѻ`,j`l�,(�����Xҙ�}HVU��&A��4.���D,��¢Dg������>P�ܽ|�<�{^����n��uy�~T�5����T�������x�����'.���/��[����W����Kx�����ϵr	�hC�D��X�u�W��p�s�U蔶��, X9�b�!Up�u`fa���Ru��ޖH� $��Ǉ��Sg�>��fĩ9,Y谱�V��u�֒9%ve��@Ԉ5P���Z]]]��ΎH� v��B�%�H�#�\�zY���CTI�P���E���l	+Y'�uttT�mDDXBX����Dxh\���<�<�����-������,Dy{kġ�;�-���6��(_898�C>��#���p�������:��^<��߇�%���\�Py]�f���O�-���`g#Uq��ޖ�U������̲/oOOu��yd~���e�r^r�Æ�W�'���d�l/��L�TIv%�9�/U�t�T���Te�-X�31#@�����M�ZbSu�S����Axd �S�������$<x�8~���x��k��������7�׹�#c�����$��������#�	V�f�wԅ!��f =OC��È �%>��M�`	M.�0��`�4��"l	P{�D;B7�z1N0Lv!>�aB�$�@'��3�R�`�����9�&%��<a��3���e{�4�&�>0��I�?�JaQ�M�0.�Yi0,+�`�)v[b`�p�ߺ��d8�'���/��x��û-N|�y��»3���pܚ [>���rlI�c{2��`P=>��"`�{�1ò1Z�.Ѝ��̥=�����;x�[�ꩃ��1��R}xu�V��I�$@ݠ����l���lI�Gy4<+���tG6���)�.C�ԡ�S�s!
��|�h�x ��8����&�N��V���K�1�wmA)�Y����T����N�h�����L�A�h�@�E�_�trЂ��P����>�\Cۙ�[xn��r�D	�)��s�Q���0�hQ�;������	����k
�Ħ�/M��<	�����3c��N����S�ڭ$6ڮ*,��ۅ�s� ��r���Yf��C;0tu
#Wg�w�8zΏ�^l��G��,k3:/�繿sD�����{/�+�n{� ���s<��n5-�a��*�hB�H�f���qFJr�s3PR^B����R[���Q��ڍ��46����	�%������SUm�FƱm�.n_���2�l߆��}O=�.��=���N4�U��(I�ш
&z��H�?7��~��;Kk�X�!ć�!�����v�}��An���P��������蕛�W�B{�*77��w�1���t�ap|
C���y��v�FSW7:�0�{��s��3����}ڼ��72���z�s��Zˠ�ɩ�XyX $;	5I��KDzg�a��6�ݜe�w���,� �X���gRź�<�x��`yXڊ�r��:,�6�]{�M���p�N�a��{	�}:3����D�hÁ.l����D5J���M�|�[����'0�Ow���<>�����;Ҥ��h+����@+F�����Y����U����Al{p�:�_��g?|}�&�<r
�	��G)�~�ƮL`��4���/��rG8�W *���!��?� T��
D��]�Nd�����P�����A0� �;Cᒿ���R *`U�Y���>���1�~��#�{��=�\�Ӂ�2��Z�v��� MF�K�&we �Mh#@��@���'����(4>��6Fß� >x������ 	��,�IIH�:��x$�� ����DH���BUDW#�,1A��
EbU�Y0P��$������8F�&	y_��MLm4�k�J��||��s��j0p��~���ޣx��c�ل�l7�e�`G����4fD��dB۲`ߑ��\�1,�3aΰ�⃃(��Cޖ ��ɅU/�,��H	�w�}��"���m��#Mș�F�m8}����w�?~�_��K��ϟ��_����<�<����:]�-3|��!��I�	E	��:~7��I����*þ�X�N���(�	��D/�uéXw��s��1.8�ɞ8�ꍣI�؛��Y�T��b��BPp=EAh)	�@[.�\;��?~/��$^���x�7����W������O�}z'����:ڍ�0`!Dc$]�]4F|
@��=h6V��b�]Jtʺec�XL�.�O�Ҿ4,c,Hƒ�x�%]P�x\�C���ݒ�$*;"��*��������P�Y/�5��|H=0��{:��6K���.+�ñbkV4EbEK4�t�`UG2���<ZⰒ�i��߄6?�F^ \�P��{?��/]��7��G΢��$�&[�ݕ!�.�)ˍEam)>��d�����/�%�
2�h�"8x��7,�i�H)����.t��|}1�._�U��AO_�Fĥ�1,�-`fO ��~Kft�p6�����D!"U8�LL�MB� ��� }]=5�̦����\m#�Q�$49�D� ���D������s��!D7l�~��Yk�� ooo��`R joo��AAAj��S�)! �
@`����z���o���p!�q4_�Gp���p���0&���dy��U��C��>� +m>�cN�K9��G��r<��D�Y��$����(HuV��d����G����ڞ �����,�ڏH�}���x-e	�0��$�``B��w"�ɹ�����G��lco��2�� T2�R�W�1�����K��3�o����[+�Po'8�X���hm]	�ęS���P���Z>�^_�kwo{�f��� )��H/�Gfqҋ���� x�x�:�
\���M�5���6�Y`ׯ�h	���F�-4��;*���ex [����e�>���; j����m�9�iZ�����Ta�)b.��a���lH��Vb�umN�OW|:2T�ӽ%�)�hO�ww���֙���o�����ΆH5F��)���g{"���4,��e��OM�G���ٗp���(騆��)���y�^�����D��w�~��j���.D�We,|��
mJG\w2Ƥ}�d)�Q2[���ʹ�,(#Z���#Wz�%@��<Ns�s��|K�*�+�w���=5��[��=ĨT�%>������
z�,K���!�ρ\Q�D���x�ۮ�ű������+�q蹓��(���;�B�K	�2d�Y�W�t	�</��;Y�l�T�e�2�#(�zy]�'�ϐ�'��2�A����͕�9��'f�}uDe=ۉ���2Fg��F݅N���{ڱ��V��1��_�F�����^C��	t��\ �D�=��=,�q���Kl� Z��;7���Xg�F�	��00ׁ��"�����bⰠ(_���}��>;�I�lpxM-�áֶn\��0}��8u�;�b����oDM]v�ك�^�{������u�QU�k�����`5�J�� ���4~���Y��+���A��ƹD���z=,$)IɈ����/��l-QTQ��=�#�Ρwh
�w���g1�}ںy�z��34�݇�����
�m},��|�������P���>~��sG���7�����2h�_�5�C�R.�����EjK2X^+�@�=����AZl�t�:�6k�k����wy}+��g��8ل�#��z�{ݏ�����i���@Ӂ~4��p�Q��cU(��A���������m�n�p'&�����D$C:�����7b���8��i\��������;���g@�_ߏ���/���0J�O=4�m���� z7T
>�7 z�P�m�3������Lh+��/���-���}�R��N$���n��Gq��
oϨ
j�D�7q��D[��/l#���U2�cϨ�&�	Z�I@%� �|ް:Y0o�G|k"	�B'��LF��"��ǈE`}4$�Yo��H�r9� ��A�����"���%8�.i�d2#�,��0�2	��WAp��%�+�Fd��J7"�<)��H�ArY0YH�+@<#�l�ZN,Bl�F��1�a������'J�<�����J�z�"���\�������{�+�
�aZ��ǖ�5���k"Ԧ9���uG��d@���a�-��"F�R�)$&����/@ �1\�-�m�@��~\x�E|E�IO�ן���}����*�൏��^Í��A��f�n�D,��dF)+u,��7'c'�9���)�8�{��p9���Ϋ��x4���y��xo����o$0"��J��u�Sa�x8�	�mq!�g�mq"�S��l�/��zb����,_L4�c�T.^܅g^���?z	o~�������G��?�������O�=݆��YFU$�{2�7�;�YФ��LĪ�<��)���\,%8e|��粑L,Lâ�,�K�bƲ^¯+K;�U,�v���W�|H���!PS��e�X��J�g	�/n��迋e��-1XBt.��ug�Y�U,�#25;���_���m��fh��M��kI�~]"6�PZ�B]x�y|����?�/����Γ���#8p�Z����T��͹H
���-�s��>":�����_��k������hCh�F䗰���
}�#����cG�����T��c����r�"T'�|ښ���$N<]aA�j���3,�*��:
�S𔬥L���WUS�H�� SP��ݴ0�a��j[��l'�-��&�@��*/1j��	(�L�~
@���3""�dAe�|J�T�S0�-d%�3�� o��ʔ
�6J���#����|P��zɎ�����J&Q�(� % ��eyLF���z]����r<9'���2��o��N9�Ux��2����~	O�G�!h��x ,�}.�9��������c�B&��e�c&�~J��ҋ�d;��e\=P��I���� ,Y�yy�x�����O>�+�>��N��UՅ(��Aզ<��oBMM>��x?��:%5���r���=�cY����0D� 6%�yqȫ�@iP��o�B�F:����j =�W���A��a����; *�N�Ʉ�~�	5��V��I�
F%*@5�:S��v����!��
�Ee(L+C�DL:4%�k>�,k�aU��8�ή�p�^U�6]�Ӄ�.B(Q�;�G>Cm����6z�a*��[��ׄ��!���
�^U�>�O}��?��?z	ŝ���QP�W�Jp��Dg,�q��G�z��4A�i|�·:�5��h�Db_!�'�T��dg=Z��S��s>$�)�N�g���s3�Y���
��"B����b"�d��"m97����ݜߵ	�X���_�t��P������k=Չ��3���NL_ن�Sc�>҇��&��oB��vt	[�5�lj!�=IH�#r����(���� ����D���d,�6m"��*�+e�[��B^V ma�w+˜��v��b�T Z{�Et�]�z�g���Q�7���c�<�7t�!T�,ss��s,�q]�Y��8��{r*��'=,�[M�5�:Y�#>%՛�P\����"���s���opG�	�!�i�gw�������g�!|����+o�yq�ی������&8;1�g�>G:��-[QX����,����LABl�ʀ��4"$1�
�;�A^�.�����!@C�A�^�ĄD���!$,n��ع/�|�j����h�}�������o���v�No�쁃8t�4v8�:01���a��ދ�.�l��Y������5!j-]�s�B�LWh,�J��0��#�$
����� �'�G;q��{0��aZb�� z�M粠�������+�7�7!ճ���6��P#v�ڋC��(��{OL����Hz­�V�z�-���� ��`�7 ;ދ�C�w���c��B���?����!���������O_���?��O_�ч��*�n���.��Ӈ0~u������ZTU��3����rw��j���BO�s��D%�����:o5���&����ݠ���n�\�v+���\'%2�jY�/�gHol����u�{��
o���B��+��:�zJ�Q���t;�GU{�^4� �g!<�%	�f\]bG�X�R[��3�!�
��� B�D��["J�EV��QH�͈B2�I�2���H�$,��M�؈deI �2M <S�d�2����3��4B3�ȟ������H+���zb�$�(A,����DbC�'
��~���C�@	�g��w����ƶoAT�\�X��6��q��܁�mLSYP�&FK�Z3`њ+BԾ/�����I�Ew:�{�`ޗ������{�^���l�BDw�.��_�F������~��O�����~�f�`�ݳ��JPH�evţ�7�M1���"�'��qOi��
�����#a�x��W��Z��M���i��^r ������9���`|�ϣ��i4�����(o����|�R�����������P�h�m�! �#1Y��3��x��{����O�!^��+��o�?��_��o~�}7.�h��e���'���c�D�t�t.�O��X:�I��5���";��E��j~iO�v����6����LĒ�$UvqZ�E��X���R�W�7�њ����p,��E�B��*�*��l#�`	���ܰ��E��s��E��X������2֔�@�&���0f�θ��a�/��:�a�M��,ffffffffff�eY�,Kffvt��6�IÜ�M�RLߜ��v��i���;�w�s,�k/���Z���B�#�Q���{��ǯ��~��~�).\>���NLύb��E�oECr�
�^E����g��k����=��v?^���%a��/���KGq��)���sx�����?�'|����q�A<t������s�~|��n$<�-aha(���8�����fFb����z�Õ����@_*J�km>U&�z�4�ƨ�e΀2l�"�F��,'��3��<�РyƧ.H� ��d�rԚ�媢�@i�[�:::���ST�媸��(oc��~��p�l)�Nd&	h� g	u�EF!�1�S&gDnA�Ía� �\�U�Zɱ8���pF���r���RXr����(d(�vF���� )/�{2v���F�eR��I���/��-��心�q���<e�
|߂'gAy�t_I5cG�є��rv�!���3��O99��ބy�WXZ�AVn��[����ӭ�<w��ݟ��;ﾌ��S���3me�΍ArJ(ERң_X����n��4����<|��{�����#)7)!p
����&��T�i�U](9�@��B�R�5���)�� U	��Z��*P�K�ȸڭn�����y�1��uP�T�~�\�V7�CT�5,��>�S��F5�0��^etʃ�]݊`��O�CC�n���X�5���К ��8w���#.}��N�Դ1
���P�&lB�	�JU~P�	�f�4�Vپh�ٍc���o<�^z5m0�{�r�5d�o�n��Q6�b�́fP���H~0|j�C�,��(�h,��ݛ-��T���p�Yǽۊ�.A�Z�r�G�Y�+�A�}R�
��@�BSg��e>�h�M�dh� ͜"(��M�:�wvXTGlXi���At�F�b-A3��)��]�;,��stT���,�#-�ޛ�br�,��DR�r?�!�N��d��H��2.i=O��<�L�]�b���%�I�M��<�p�*��щ,���~�^P���ݨ=�)2�<�!X8����D/	��g��0,�	Q���[ �<Fe��"�� et�2gH.L6��S]/�n�F��P�Q���"�tP\Q���1TT#--�i���ACs#��wcyu������GIi�����<ffw����]���i�mC�::@���~S���ANnr2S������(�D� $�>���2W���|���t�e�v���w�h�_ �c����h�Ϡ� x�� 9+�]���PQۄ��VQ���}PT��G�0!~`��`��^X���Qw��>�Xً)Z��gE��in�W0��,-�i�eMe�+o��[�z��P�P�G����К���4_��9��g�����]Z{DR�6	��|���P΀��o@�J�v׉(t��:WGѴ$(wDĽ�&S�3w�3��U��~Kͻ�0��� �~w��?��������Cs"��?���]X}�0.=�~�,{�Q�|�V��`��e,ݿ��/�Ğ'V0~ic�>#��o *�v���7����;�vlJ���b�X�=@t�k~�	P���{gж�4�v\�*��DZ�ǽ��cS������:igC���}��9��,��nK�s5\�zrU�f:�v����U�LD���k�@tu("	o��!��fLݤ�c��(�T�����=��QAA��(��Y�?��Dh�-	D<�3�$@�3�PW��g�3������D* �28)��	>��BA �P�Z�Gz=A11�I��,
:EB6�6�Q�li0�k�L�5O�B/D�{�p��C��x���X\��
�U�tb������@h�B�(T Լ1	&M�����DC�*��Сk��J(i�%|���?fݙ0oN�>
��}Q4ۊ�/^�x���3|���������7����]���ѻ܈�b��Y ����a�h�De�/*�l�f�Y�^os\q�#�v��k����J�=ލ�����pg�G��9���0|�Ob��1M?�p�/�}��?|��o���E�/�u��J��>!��X/�l��,q3�g���Yc��h�TG��9��㗯=Fe�O��o�Ňo��W^xo��~�����������H����SaMa0��ٸ�йn ���!Bi_��&g;�389�i�7���=�{�M�X��{	��RAfC]6��a��%�a]��E�b]�+6�{(��-��b$�ì���}O��|��Q!`] M9,�.��#��7(ƻA=�:��0H�iZ�+���q������7���7^�^��0��1�c
;���g�em�Ȯ/@ryRK������(�^š����%�%̎�Wc~���+��sg�ũ�����׿����s���?������9GkK�l�,`ac
{s�(!���60"��r���R�sp�<\w>�q�[5pgBOn���%8
�ji�r��1��H�)i;J�UT��� ��>4�8���P��`<2(��L�l2>###E�[�)g<����)�+O�hF�$+h%���z�C��1
�*-C���P�����ؗQ��1�}"�H��R>#����CF��<�E��}���|}��:i֔���VZ:O�Ԋj�t�������)�vJ���zF*c�������f��K�S����Ѳ8_��n�'#X���ـ����o҆�z��ˊ`�:��^�𣂧�=g��[ ��O��7_�K�<�W^{?}�1\�z�,����i��􄛧5\���n	[��8����
��aQ��<l����p/D� :1Q	Q��ߔ��P^��BU�ր
�s4�M��k%�"T��*���,�J8wF$A(g>�P�~r�\�!����@��\��F�,7I��|oh�C9����R[�?
_h�3N��uZAХ�A}$L�fE�ؑ��8��e���iK ub�����5���ЫYO�2ol-�B�Tj�^D��czFz�Ģc�0�>s	��~���h�9��`&zJ J��h[l&�n�k�N�z���&·.���1�8����\Jv6k	e?���H�q7	�Y�\��YЌ9�)w�@���}�z�͘)�i;O������P��
�{��j��GP6W��ڿ#a��u�����:�me�d)e�P�P���<6l���!r�м҉��j$нr�^?��T#W��b�R�|*�"�p�>��V]���*@�d����N �mi�PF�H�$h�a�>CǙ�A��
���čy�\ ���b͉��#�r����6���������)^��ȥЖ�T�#�J�)�yr�'�<EgDk��!zM�l5��黮�{�7`���IU[�vf(�(��� ��ˑ�����F�M�blr����Ҟef/
�K�؞<�JQq9��[���Iϡ����fTTUcxt��va~a;�F�����W�������`?��@���@__X�}GKM��p%tr�ӛ �0��{LrB"��z��#&6��O?_8������Ξ��E�5�smh
3�{�3h���	t����M]��Y�����t�|��PΎ8~󻗑��#�Wj�I����
|�*n�&���W�^�����������@\[
2F
DС�f�x�nUp�Qs�]T�0��|g�S�>5�n* �Z/��e�û���U��E�2Awg��g�JJf��E�/�� Z�G�	Q�r3��J���]����3�"|n{x�.|�=���g�rt���g���O@��~��a��p� :qn�@�.-b����F1wq	{>��/ݏg�7^{'n��e�"�rP����q	@G/�c��>�=���Q�_Aߕa�\Bׅ�!�@Ȱ�3>�������;;�P�v�(�#Y�5h�Rx2�迪��!鱖�o�t�|�}�U�P܉Di��[�9�=�����I�Q(������@*�w�y�#a�σ����m������A}g��O�('9��5iG�J5r&�f?��dU|m��O���E�c+#���	��U!����,�A�/���^�. $��������B|a���T�d��zP�2�T��P��ˠ�}	���l�b:7�
I.HN�p�p��A�!��S����"���V c��C�
��q��<����/c�� r��B�4Iq��E�''|�uFdLt��(�A>�Jt\��Ph�E��/ڝq�h��Ak2���ܔ���"Tʹ��cg�������~���x�������p��fQ�)-�H�@	���6Mt���q�F��6�{Zષ-��Ƴ/z��u?;���O\�i�;>rÇ�n�8�Ez�}�(�-o|@�I�?�$|~��_%K"��i���O�]�Q�3>
qٷ8C�k�'|lq����b��HA"^=4�����W���/�ķ���_�����^z
-+sp�ρL*�B�֓��dlN$������(��t-7�r5�p��cv�q;)�B��.�jC��
{ύ�=\���i>�������ۇ)��@1��{�>s�~;�TxXF��]�ڿe��(Y����d{����vS�]���������B���\��x8%�����^x/}�&�'x?z�<v�!<��C8s�V�,�����߳M�_�Z���l$��!��"?Y�q���6l̕�b�/']��� �>���bLN`iy�ϝ'�������?� _|��}�M�?}�
�PWS���5A��.v�q��%��):�ч���p-�ʄ1=1����E� 5��oU���p+�^���e)@�����9�P,gP�*/C����Z!�K�aH2,}||D[P�wuu����j��}��W��m�k���(]"�I�g\2*�7FP�ՔB�q(i�)�N�k�\U��ŀ�y>���+z���������Q�׍�Ï��c�90�Z,���L�H[	Dy_��~|.��"��� %@ڿ'������S������ʜ�e�2��<�`���y�:������q����(g¹�-g@���>��aF���� ��`��������/>�'�zg�����k�,&g��^���@�Fz��Ò�wư'|Z9�����J��f- ���D�uE`�'���� D�!&)����
p��*C�P�*P�ׁ!T��*��P$�ru\E3��6��o���jQ�6��M�(W��L(g?�	�Z���"�j%9��~jf��̣!T3��y�P/��
��C��j�<�Р�:!����0檵MѰi��m{�Zba���v'���H�ik��"��. �B�y�|*T�s���[�"/h�{{��c���{�a<��M��yՓ�M�Q�7��=�%����C&�
r!VP�p.Gps:���]O ��wm��(u��;�?_��I��l)��)��9WF�,á�8��E�aP8�&��P�����kF��6�TЮ[m���8��)�ABg2�KC����L/8p�ً>?[(Zm�����CNw=T��bD���"6��STNV�s_�	f\E8��!�QL�̞)�m+�yI'E9�t�S�LF�$��/gcy?���Ѥ�L�k�ȢrD�T�)^��o�O�(����o�)���e|r5܆�"�K �6�穬}a='F@��!g;E��S��n�|J��-Gz�6X �PGl6؊͚2P��
]cM�ۚ <&qɱ��ۂ�<�a`���	7�����A}cE�[QG��̦�=�ťU����;������kF�� �m����a�	}�Tnno M��@tx0�(b#�	?��r��j����CNF�󆽕�}|���475abbY9����t?�p����>t?�&��cq� ����0<��s�8t�,�7���n�w
|�;v�=�S<�T6;���i;w�/]A~E%l\=`H�0nc���
9�-�Q��f��W� �-0p�Cdq$�;2D4m8-G��{~���������Ҕ{�m8�C擫�����Zf����<�*����~��G[E5���h�ߊ�K�Xzp�G&E�����Չ����Q9�/o��(�و�=�b(�ڽm��K�#��a���Ѷ�]h<@��[mF�J+��v�{� �c���UwVd@��w �������%Ї�ʋ�E���x'=��KK�޿��9���� ����T�gA���Bq'9|���F���ø3)��q(�-~P0�?�OBi��|��qy�P�|r�d����N�>rPiV��~����?����4��� ���eAH.EREa��1���pD�(�h ��_?�?���!��Fh�&0rF2��J M*�A"�2� ����|Bc�;�aT�.��J��w§��\�F�"Ȧ�JS���H�HI�pEJEgC=O�퉸B$UGµ  ���OqCvG6V�l�B�	\p;�� �,v�v0��-���^~0�+caZ���G@�*:UQФ�U��Xh�E¤?VC9�� 5z�=0N�����bL����s���Sx��#���^<��^,�En[�+C�\���䡹:�tざ��2Ñ0<��W2"�ZB ^�����x'F��|/�?����.�����w�S��x2�O����pw<��N����O���"��f�/~Ι�5�~�/c�	�.RO|N�>�����i��^��1�+�1KM�9bgy:��9���}	��/��o�����a�̋O�$=?	���t��U�R��'��=\�6	��	��(�m
�:�)<��=����pl���f��ݛ���`d�L����?�
����x���⭿���~��C����x��?��}~������g�+��7|��?����Oh�/�w|��������3�}�M�������_�᫧���><��x�w��W��7��������������g��G���C��1�6hy{2�r�X�J��$$e�#=3i)!r���b	�yt�J�bPEP�l���H������p�ƃx�9�;_}�~�>���s\�|N�
uU��z����QѮ�q�ce�@��xh5��&�9}��@���TY5Fc�A*i�)��+ J`�)gKE�E��S�UMI{P^檷�P��˝�b��
��� &&�V�Nƥ����;,b��:ΐrv�!��y;C�����P򄳙f�LiUV^�q[oOO���dAȄrf�����'2�|l����>T�b�2Z�C^f�qF������?�ÔV�e����{�T�`˘�y��)��D~oF=�W��fb��`�G@���u܉���Z�����p�[����v��v���ցA���P��䎆��D��O��2b���� 1�(�5jgg�-2���%���}��y�5B�8s�0ك��I�u��>��������=\<�a�F��}���=s2�5����$���!^��'��#*>�)Q����	�,��a�5��9�A�Q�κP�&x��@އj
5B�V�� ���O�z2<��AEp6�@$2��N���|���lwhQh�H�A�V�	�b�[ �"T
PMz��@��`�	S
F�U[,[i���$XS�w�ø5M�����P��"�S������N���B�=R\жo��~�1��*j&�a��X7e^�\pO�9��@&؂p�)��"�6� �Up@�$ -Zl�pE\h�M	x)���D!!�@7]*"�"���U(��F�j;�N��� ��|����xD�ESD����%{�Yl���,dL�`���n�V�-P0�EI(�o�*�K�\��P�R�[�*'j�A -�V���b�c1A���Ɣ�9](ڔr�|^G�d�f149�9A��t_ΆJ����\�w$K@5a4]d@KWj��)���ð4R����r泆���d�ta�P;tT��ñ0@y��}T���������)]�;ǝ�!�?&~�آ��z�P�����놶�V4��#�� Z�O��BO_7�G���َ��F�eZ���D�dh�WԠ���b�EUu#�:�L��I�u��ߎ���clb��u(�(������[�gXb�����`�ҽ�{�5�7DAv.vm�!��{-�[�=(<�UU�=jZF:|�E�3)=��x����72J1�م=ض�OdA��-a��Ӹ��T{F@sja�=���|Jĥ�ɋ�Du\nʝ1T�#c`jo'z{�0Ԃ��VlR،M�[�Aa#6�n���B����C��.��s��7�<�y�������u���[�x�� J���#��5S������x�5�jo�W�0se�?~c'�й:����]t��]"*hx΀V.K�Jт��&Qu�e� hA�f�Q�m�ӂ�}�����m@�ol�ăsb���1@/��^�U��>���z� z���t��e��Q,�X���i�<0���� @�w���o��w�|;<�! z��'������`���Up�|.���^���6��}�^po���T˵|�Y����OD
��Y��Fc0��ÑV�$΂ruܺD�C�����
BPu0��V�HgL!ݨr}�ツ��!�ȟ���d24�ИK�� �J�鎄�f�J uEcs��T`�OuDB�#)���L MNu����<��H
�(�:�9��Lv�[�?����6��1\�����ė���
&v��0��Nw� ��PWDð2
F5�0oNUq�a�����g¡/�-Y0�
�_m���Wn��·�}/<s�N�az�mÙH���	�Ua�'̖��� �E��hv��~7S\r��R��VN^K�Q^x.�?%D>j��!�x<�{Y� {܌póI�x�06�ዞJ|=T�_���������W��r|�Q�����Ve^ʍ�O��4a�i���"��"!��� |�%�~J��O#=�I�>�����x��
��1���ڛ���gG����O���g����;�b��2�g�����5��5��M��X��Ul���й�!��I���Ox\�?���u����Qq]E�%,j�q�˷�1@p~A���὿}�7��%^���b������x��_��?��|����������x�᭯?������~o|�6����$P��_���y�a��|W�]�C]��ׯ��G��}�\��kg�g�.�����u�H"|Fe� *%R���D���Pz�#'=���(JAME6z{��m~�� �>���}O��<^|�5���G���p��i�s�>m5�������F0�0����m>9� ��Z�SX�8�P3Bg+���&W��	PJ0��8�Uk`��깼c�;�	FB\� ����r�S
P΀J;"�*�~~~��-W��ඡL�r�2R�Ps4;)�܇Q'�2ؤ�� @	�8���3\@���&Ï���c1:9��z����\�8��ǔ�-�2��?i�S�:~/Iv�u�Zb=����yJ3�R�r[P�+.����YS��u�RW7qL>6W���� U�	e܊��������QqulEEQ������pqs����;�U~L���ͼ�2�qO�|��;���`���O����
����Hx�������PK'���v���lkK�z�=���� � 7��""&�q�HL�F^!3�E{Q-Su���0-��p6���!����P���Ԃ��f}+��YOi�Oi�Oihs�B'���=^��z�l����n�'�院���/hzC��*��e?	��Oz�iW�@�6�u�b�Scz��DK�ٙ(�gO2,{�`����73@�<��O�j:~S(�ڣ�x��K"P���i�?��<�s*��r=;Ga���xw�g�B#���.�I��@�A�3��O��$�g@�
ndw&a��;�P�؄��*��n9�9Q�th6�r�W�P�܊��(�V���Z�"�!EA�|t�	�_�[�Ϊ����F��`�8�i(9Y���@�B�@����ץy�-�ז���,�͔�l�H��<��P<\�Fz�� }��]�%o�X�������%|��I	J�۳&(n�fpft<�R��󗳡�4y"E���c��]C��A1�g�	��Zܪcm" Ah��gG1ruC��0x~J �3��G�\FДb��)�~+2����;/Atk
���QcT�����cD�Gb瞝�Gem���Չށ^445�� ���-z����A}Cjj	�u��o�i�E5�����a���:s�/^YP��('/�9��ml=�b#("��+ ���
owO�н1<8%�(�/����(�$'#))	����짿��~ڻ8���GN���"�zz12�M�svaC������VőS�Dv�3��;vR,bfq'�<�s׮�Щ�b����Sy0��+�з4������QaT� �	��2��#�ʎ�i����x�o���:/��������q�Ҷ���o%e��TZ햷I��@֨>چʃM�$���i�,�Г�0yf�hZ��[T��aX
�j@���P<_���zT�n��Upy��z�=Mh�׊�C䞃��KH]�G�;yx Ë-w�vn���({�mDo�� ���N,�Gb*o���9�k/? ɀrP��%�vߑ�N��Oɀ��1D��B�'���- �foe/i^dBy��h�yg܆��i�1�y�P�1��W�e|r�O�]�蔞�< �C KEzo<Қ��Z��� d@3JC�^����PD<c�#]���P�:������6���-"�#.�����3@�~�MgR�7�r��n��rA�3a����g��ӝD$g03\�‸tZ瀄4$rB�i�L7DS��k�����P8���*�M 4�=��Gq�~KG�Mbt������C@}�����4*����,RT�ի��Vi4)t���_��hض���5��O��(\y�i�
���_��^��<wO?�;����3F@��j#Qِ���0y���D�:��f�s��x��7�P������^��a�󞆸�g�+���m�
"�~s���o���>|�{ �^��=��,�K#�n����V��S���c�'��K���!|�W�׫�p3=��]p#�φ��|�L���Ǆߏ��A�=��ó>fx��{̕1a��173���W�?��7���_�K�o����O��W�urX�*�)u�`c[8~B�\�=��J�����ý5��T���^X�����A6��;��s�!f���Ɖ����U4�ߞ3R���r$u#�-����n�Fdc"2ٔ�HZ�K�_E����W�����P�T�+�^&���G��?~�K��y��/	�^�r1@�H��C��ߎ��T7U �4�9�MCX|"cC���̌dde$Q �T/�KFI~2��s02ҍ�}K8q�ރ�����_�O_z����׿�����r��������%��L*�m�agoS3�de6CS]��i(�'���P �aɐ�v��MF'�g�HzV���j�7Q� �L�d��FG#'3�B^��d|r擧�K%gA��L)W��j���/s����}����>W�*��σ���B�3��N�3�\��Q���YG>>7ITҮ�;⿛1�M������]�[�������d�:���⌨4[�ד���x��|�"�I׎���M���C"~ޟ1���������%���9#��������܃1���Ͱ��U�s��o����5nL�TRU�V9�e|�9����.�����AqI>�}�M���x�gO�ͷ_�O>�c'�baqBT�mh-AvA'��p#�:y����F6�0�5��}.pp��;A��~.��B�361)�q�i(��v�����*�j�A�T��:Pu%dyB��{Peh�%T�-D�S�.cS��S2$�r%�W�ݧn�+t3�$ %|�0>9�9�S��R�8ת�r��C��k�N��h�����%��Q",;�a�K(�Ӷ/6V��0�N�q7͈�nKT��(�P���p��=���ӳ�ۧ6��_����{O���W���X7h&�C#ӛ�7[��Z磏�x��?���D�[��84&#�=1�9�2.�#{��+P��e��w��'gWZ��ۄ���.@Tc,�
|��_C(�*A�LF�2�b�	��[ k��4�`*E�P��+�E𼂶d���<�5� ��[T6a����V�[�B�Z�.z�H�F�Hwu�t[=r'ː>ZH�,�̟%pNK�Y��PZ�Y�g�t!�f�	�y��M���\�ͤ崑l�g	��L����(g@�'\���&�(�;��2W+��H'�OS� :ryFd@{O���� zO�	\2@�"NH�fi8�%��O�z��G@�R��n��.T[6����������"���-M���!WFQ�X�����l� d���N��\ն��ʘ϶��
|NN�aj�_?�CGc��E�W�����Y鈋�ð�E�#&�~����`��������0$%$���1t��,�����GjF:C�l/[�!���r��˻006���y,�>�]{�`rv	��1�}7������>y��ۂ�o�YOn�ə���{����EV������6t�1���}��
���߈�[���FX��#�9�P��[��
=��wu�>�Qh�`�V�*��<%�����:�P���h��'W�e�V�oðL^���G��|{���h�R��%�� ���Z���?��@	�5+�h�,�F4Ҵ�`Zu������~���Mt��%����W��O:e�_�����~e<z�_}H��unz��ڀ.?�c�������@)8��h�cN ��~ݝ�?(�N��EF�J����pp{�nڏ���p��G��gCy�F�5�j�I M�Br}(R��YLhhq0R	��e�H���=�EԄ"��a��� �����@h J��XD% �Q$"�  I�~"�
%f{4�,���4��ጸ4GĦ2i>1��S��n��4;�f��TG)m#�Ff����ވ% ;.�c���ܮ|�>>��oƹ����>���!�&¡6	���PN�Z�/J$�@�	��Ԭ)�
�0oI�U]"�*�aDp1OCVo~��[b����.������~�^�GC["3m��D�nYt�����Z�vX���!;=\u6��f��D���Y-�T�1-\�r��x�+���᝶l�ޜ��+cq%��ݰf��~f�#��hwxZ`�
���]���	#|q_N/��s��x��7����n�u�/Ue�Ɍ0<��c��n�;>�t��!�x/�o���Ec<�k����p�QS���B瑆J<y� >~�e����?��/���=�(zW'�R�u�z�T]�X�,�yo-��N��u������PA+��-��x���x
��}X|�A����0rdi-�0�p�|�1dC(żB���rl7�\�!�h�|�!�`��6��T��-^� sQ�^ ��̑\��z�����W_����w��>���8v�Oǅ�gp��)���#�`߾]�>O���n* ԣ�"���I&|�D�!0& aq�H t����$#16�Q��H�FiajK011���Vq��Y����x��7����/���������W_��
�*
����9Aʆ jgM��,AEI[ee��� ����	W<�*��MI�B1ϐ�L(��&�SS��3��/F��*��BV�J����~r�I��SF(g49�Li�C��|˙R^���6F���#g�\�VRu�Z@�q�!���H>W�r�v^���j��=䪱�O)Dw\���π�GҞ�P����*#�����׆;`RVT׍χۦr�YF&�¯����0F��lRB��Eھ�ύ�����q�b	Z%�O��,����6�����%�$�����aF�����nP�R�2���m@�gd���mCy�Pn���͛�#-=	����ݯ��_}�/��7��/c~a\T��m,@ZNB����g���,	���z0 ��:���˕�3������	�@p�?b�"�����������h�D�%+QW�U��5��>�7���.���T��v�������47h�8���\�VWT���T�ͥ)='t	��M��hWC�*:4�K�j��0�E��-���p̂�`6\�s�<�)�z��ǉ̧m��a3�B�Iw�	�m���궍�P��AT��茅^CL�=l��P�܃'>xO�tן~ �Kt� ��N�FE�?�3<%c��Y£2����oH6� �5�H�aː2V���\���!��;��mV����vi�0����9'y���B�Zu7`��z1�b@�4$x�m�V�-��و��P���� Ume�h@�(���D�
PА���dT���flPވ-�2P&��8������(�Bݎ6��ա`��Eȝ*E���%�f$s�
QL-�+��K�W��|z����S�?� ���8<�A���S9�ICɞ�^C��q�jz\�.�6�2|��6Be�Ȁ2@Gg&�w�~f	������8�ٿV%w������*xA�J�4d���
-]u��z���#�èm�CQY)�jk�?8�ΞNT�T���[m@�+�h���}�����4��;�l��)z��ݶ�啽��9�N�����Ņ()/��y2�cGe��x�$Ĉ*�I��\�%�F"���C��EŠ����H$�vvu�yԢ��Z 4)��oq1�v��YR<n��i|��/q���]X���CXZ9J�+b~��#8|�,N]��=�ctv#3��������|𐘮>���O��g�t.���0s����6�4��II����c��0t�EhU���P�̩b*�c��>�f2W�e�r�Z
P�b+|p��J��Z����� e���N�� ��@��b��8��-����B��~[��	y�H� �h[J�P��	��L%�R0<�%�@@w����;'�Y�����7@����0����s��.l{�.�c�@:N@�6��ˤ�3Ch������c���0���Ә>K=�s��:�]܅����+���� �>�c���K�M�wݷ'�0���*&�La�>:�x� �1L ����Q\!@�#\u����A��[�Ý�0�x��;q�����O������n�nm�s�=�����[�i4s�k�������/ڏ��H��-�~�V�R����tm�����\Ndo��rZ�/K�焎������F�?��]�ov�K��H?�����(�ӻE7�_��a�[�}��\;�tl1�=�O7]���:�g!�9��Ȅ2�b�?���E�2�8)�AH��T�S�J0Z�HBjtY͇ ��c�\�5�4��LA���k2M�i�X��|_B����9^"�r=Ű*�Yn�&PD�� :�	�Tx��il�3���`G79��I���$9".�q�J0uGt�b�y�QWz/�4Wx4�r���6<��9<q�(V�#�.^T 	��A�@;�`W	������<z��0!�z�s�6-i�&�X�G�(��g��/>�W�
�|�6�{�~������b��"����bW��x#+�Y~&�5SE==|&�����{����H�m���B�MԱ�H����厷ۋ���]�G�cp:�Kv�X��ڴ��td1�/�Y*��(c����(b^G	�T(X4Ҥu���VĤ���m��X�"��Y�z�>l-�'�}��|'ޮMǍ8<��c=�L�����K�.���=���M7k<�a�snX��A���\��,a�>��?y����G�%��~�*�r�qvPh��=5�XW�u5^����Jo�[�u�θ7�	F�(�0���Qsa�'��I��l�9dB͡[��p��D��9
f��T`���M0��ѯ��eU ���3k��IC$t*�`���R8�$Ø>s��@��K��O?�_|��}�)��٧��c��҅�8}�\�ޕ�X^ڎ������� =�+QP���8D%�Q!=�~bl�`��E 6�~�HK�Fr\R��Q^����*tw�be�zx?�Ǟy/��2~�ͯ��}����o��oŕK$PW�G��'<�aog!������6}��S��С��*�F8��i�'`�AM�
���Mm=¦�����e}]}�����E�s����K[�����E����A�D�O=B����@È��	�\Յ�iI�bXr���b�*����C�H��J;*b��q�}#O�s">�-Ñ^�aʠ�m�1�ET�%t2~���~�C,�=�Ж�� ��1�����5ԡɘV��!��Z�k-M�`efA�r6��������:����:|�Z1p�ܮӍޛq˰��)Wcc��g�ׅ�v��^F.�����0����a��?h;�_��S���Iy<>!�������.�.���&x���HYUY������k��(�c�"��a���w�w��~��x���x𑫸|�4�/N����5�HH�O������<��a�d]����i�N����>f_G���+����@XL��P
^vr���>�ԡ`����:P�dx�C%�
j��"��-�C�x;�q�PO��r�4�y���!:�� ���@#�Y�f�!�"��z%�0��i}L�BaL�WD��H�o�B��0��a�g� A���5���T�M��i8��	�pN��T&\�Ra��^��Dì7Z�P���R�t� ���.߈����~��덟�č�Ǚ�/�wa.�AЉr�n�7�9���z���߯K�:�ӯ1	�-ЦD��HSד�ľl�t�#�/�p�l�x�6�(��M��b#�5�0�0\���z�
t��o�f�MآJ�T�y2ت&K�r4��子W����CQFL�l݄ͷb#6�m$ l��6�\�.z0�N�ҽ�ޓ���z��ՠx��\Ux,y�N&��Z��ⓦR|r���f��!k-���O^/��r&�2�%�pwN���� �.P����@�:N���!�z����VkEgDc��a���]�ʎ��>Ee�3#�w��T�<BX!D4�r�1:�1Zw�ʬ�����A����*�L�i�	Scxxbpbg�\���$�����M�Hg'J�ʐ��/�YQU������cxdc����&���ԁ��z��srj�O���;>5I��"95	�񈋏AfF
�*.���&�@�IHMJ���0v�\FNf.��9����Ʊ#�1<4���,�GF >)�P[���w^��ty��oa��2v�^���2�m_���"��>��'�^���nt��c|~G�^�ν1C�v��ƶ�����(�chz�))p�񄵧t,����El����nQ�%*��j�E��ț(Eӡn,>�۟Z%���`+��\6�2�ݢ��q{Q16(���d$ΞVjA�f��j��v>���gѳo\Tí�с���(��ERw�GKP����j��v�	u���x�΅��4�`�6�kC}o�t�s����0���Ư"}�������I ]�<!t���~hN t�
�C�&��^t��1���?��3��9��_݅�I��}�C�?�>}7߹����"�a���ǖE�;!�:����ϡ�c��WF	�?h��
��s�r���l��炇����ւ3���l]���'��2��*-}y��V��h�-ڎ�8:N�S��� J!�%���U���_h����4�w(�N{�hZ(�_����z�2@ �"���w��~t�t.mG;���+ �{�n�4m\�G�H&��W��RBb������B(w"T���0I2���W��%t�rƓ�GӄbB(T��H �
c9�1�P��\��'b��Tp���lT*��"&�1�NP'68����G�$R��)���xY
*����|�Qԓ���������reK+(nMD@�|*Bܞ���\B=�aN��Ր�&�*��҃ު!	���p�M�V�KR��[��/�~�ۏ�������p��8��H��Gr�;b�ꮍBc��*�41���mT�ݡ��]�z�f8�k`��%ND��Bj(��͚\Ϗ�N/s��`�@sF�X4��nK]��g��#�0;Fq��'�}��P/���S��D{M	�F�i��},�a�-��m�����Fs>������xV����@;\�ó1�x6��y;�IO<��'�\p����5�c�sa��P5�z�$���C����?����Q�+��A��S[Cp/���*��
/����O��qO�+�8c]�>�jB��ڊH*��7�����e�b�D*�%����u��y^o5�ˁT�Ҽ.aV�!ڄRmn�;��mU��L�N^��0~?^��M���{��書��C�v�Ο=�#��bi�<�g�156���.ttԣ��YV���L��������P�y�/�A�
�Dt�/����F ���ZZ�E �F_o'=�w�̥�x��'���/��7�����������׿���6��iAMU�^�pw���5Yb*�e��1���T���$OUYG�.2�s�Ƅ+n���}r�I��O�>ME�ʴ����CK�ۈ�8ywP$Y�K�Óp�P�$r�P�Zr�X���A����|}���0>y^�D^� �O:o)@y�۔rHۍr�]�۳��ZF,wf���*�<��J���zz�H]�$W�5!D�������Ҥy=�^֒�Yҹ1@-M��z��*j�KmuQG[{��{���N �3��F�Nr&��9xY�yg+����%g���q�����m�l.��a*9&�#J׊�*���:��\�L)��� e`ZX[�v����1@�eŔ��r�a����Fvu¦-	������_~�){�a<��\�r�
���DE}>��>anp���G����f�!��}�ԑ��͊
�6��q�=���������CpL "�����P�вw�7L�j�:P�׃��ܩ��ee?�:�l�l�hkѳ�&��(=thz��b��${��8B;�Z��"o����2���!0��YM0,���0��M[4\R�ҟ���7����Oz�BۼƲ�3���LxL��u,�ÉpJ���#�pO��4�o��/�9�L�zm 4j����m�Ns(�j�Q�-z�q��w��c/?��O܇����L�^�+s��D�1�7ȥ8@� ���Ϫh���mN�WcZё���L�n�Um8s[��$h��5�R���"d�B�V[� o)y3�	�҈
�:[�Qy#�7B�P�D��H�T"p*m�U���<d�n���"Gx����شu���mO�_�&���0�=9('���V�d[����d� #Ò�)�&#��6�2B%Y�5��kn��ϡ���l!��3�(X*A��&���2E�.4�%|�jCՉfT'@�5��@=ꏵ����#�g�q��Ie��T.=9H�D;��:�\y�� ڎFh����z΍�Li�l��Ys�da`�goG��bi��=~��T^#������K@�������gQI�^ebj�v/crzݽ}��o�}ZPQY���"tv�bhdTTۭ�����h~a6Y����HEbB,���G��LKG~na49Yy()*GH`8�2Q�_��dn;����tRy0&y�������ܼ��7ԍ�'U?�  ��IDATcrv��=��lێ�������VV����cv�
tS;v�������	�-�b��Q1?�������s�1�s���;_7ؚCMO�*��ST�fyl��(���7��В�r䏕��P�܋mO�2� ���Oe�6*K����Zn�ե�D�`��0@�"�5�6�c�&�p;@��M�se���OQ4U���ld�x�
;��+5+��G�$�6JJSQw�͝�4]n� t�b��d`r�.37�c�q�����zh�`J���=gGė��~�_ ��!���O }��G���ϊ^p��.���}�X~pY���i�� (ge���	|<<%����]��n
�r�Vdj	u�E���9��]��@�ܭ����;�����?,-t��t�m������(�ϔV��=$�$`�]Γw(g9��I2�W� �G����;;��~��YT@���p\cҏI�� 4j-�)��Y���@Ds���-D�����@s�p�Шt($��T��%�F';8M�(��;DP�#2�0��D ��$�!2��y~����J��<�q��� ��Y���DV���·1~���zho�����C�{,*��_]
��x�Ѓ�Y�%x�˷��o�}�<���g0�����H)p-1>#l�g��&t�`HK��Q��i`�L#�X�ăEqx��7*Sp$����h�ބn�-3QƂ����u��Q*��7�i'K�w��gk\p��E{K\�8ko��vf8ek��v�8�`����8jg�}z�m��yE��mƬ�2X��h�ޞ��������%m4p�� g��,� �qg[<��nv����EC�ƽh�P��b|�����~�gn܇��i�,�ù"��� W��� ���ĺ2h�'6@�@���c]�%4k���	P��,X6Fx:���=)���Q'��
��i�`�2>���`AH]Z����(�pf��p�e��-F%��,ƎK���O�/����zO<v=p�Μġ+X����P/z��\W���|Q��8?�Y�HJGd�B��H��#���p�.�tED�����$(a�(7-5����y�;| �>�^z�U|��'������g���?��gJY55�)l,	IV&��%�Y���P*�
PP�#�*X�$DB�1W���k%A��c��Ked2R9é�ĝI��M�xgA5�4�A����s�EUR� ���2�G\e����S�/�"W���bJ��26��q����hH�cx�<�����NT��'��)ݟ���*�_� 5�׃��9�
Vf���,��ƒ�:�}���%���� V@����|��%2���j��9<]	.n�����<9��Ud��y���ڰ���$�i+���v��Ɠ_+�Wy�:I�b���J��Ն9x;��=��w���m�y�O�Ŝ�9�=�2B�t4amk''�y��1A��mAzV~����7�� �!n>}C ���X=���k)AF~<#=��� g����r�60�'�;��J ���'�:���	!���m�cS��%��D�����V�P3ӄ
!T�A��Pech�[A7�F�.0�q���M�<`F�z�TwQ�֡4�2��x7%��=���)�D�D��J��P��HZ�D��R�N�#�ǻ�a���N qg-���!�p
��"�@;moB��N�8J��G��\z&�
Z�����V�����YL�v�E��a8�}J��c���Nk8t:"�Q�lGȅ�d�?��y<���x��0}`��"���,�5��C)�����Ht�[y$»s�ӔHs<��>ߗ��<t���<��*�U�|w���� ��!P�ֆ���](ՠf�
Uk�X�`���+��B��+l���I�p)�[���!�U��e6�s܁O)@u���P;8�zç8����Y�E��ș,m89{��g��O�~+ z��� ʯ�)W���E>���>o�g�t� h��t\���	@�ϴ���Yq��G���.���6�PYz�>nZ7.j6�r=!��5E���nR�6�A��^*�`���/mC�\�#l�Qc��e�W_g4w5c���zP�m<���G�lj"�4�9vRy��961���.�aa�~�S3hjn ��-@Mm��0<B��WTV�����Y ����Qn6�S���EϠXBh�fg�weE�HMNAJb
2Ҳ���'�&d����UTV̠뙕���hmj����	M=-�%�cf�4�\<��gO�=� y���\���FǷ���m�T�ډ�{�cb�.�KF��}��?I�ZX�O�Ǳ�W���`���,)�[���;L��i�E55��}o��� (��쁚�Z��@K�y���+`;�t��(}NT���Q{���v�)G��.�Qټ���c��iE��&T�mcx���m9>���h�=���ԯ4�+G ����e;jQ-���G��F4�oA�����#"�ߴ�mC�r3�v�`pOF�;$ �|`Vm����<@9����-��P���趙��_R��n �9?��5��_څ�T�}���������7n��#G���N츸�=���W�a��^�_����iI'D��'� ���!��.�J* J��*��ۃ�Iaz+h=��ԝ�J�[��������8��YOΆJ{���(ò��G�ɵ�w ���;;���3�2q���n �$�r5b�2@��a���ИR
��KM��,�'��#��"Ϗ�1�~�P���?hT&!�����t7��4:� ��(��J�i�p(#T
�hhD�'"�"JC�Y( ������h�������S��k�EDE|+��Q��vf r�)��>\��8�ú"N�Ip �Zd �1s����K���^�k�\és3��CAM�,}��OW�1���g��6Bf���Ԕ0���>MEZVB����е/�'�p*=cܰ�c�iG=��cHW;,��bg�CN�8D�<�H�t� \�$d����yB�y{+\�%(rB�ٙ�,�9�３N�묍p�B�,p�R+���n��i%L[�������;�Ux�<	+~����s�j��W�1-�3��ec=\6��YM7��2�Ws#jp��_<}���,^{�)|���~��� ޔl�rBh�6�{��/��O�.�!H��E�8R!Ҥ%�abj՝��+�mQ"�:cBy���g�Ƌu��T�눆fc����P��n�*wq���C�x#Ǝ.b߹#ؽ��]�;p��1�5#�Z���� z��T]���lg%#/5���QH�
BD�B<��?o'�x9��������;41!)	�HM� mo����0v-`��Ckc���O�����7���������&�3����BH���WݔԜ j�@	Jʊ"kȸc����s{G���1���2B9�)����M)�K3��Q��B]���EǓ�U��UE�����']�h��G��&CQ��d �2wN�c�J;)b,�>�K^�Uk��.o���M>���Ҭ�4�����gNMyjlks3�B9�	�6ְ���2C����%e����ٞ
�N���֥С�[�k���rد��D�!��� �br���`�PSï��z\�����6��:i{[����dxJ�)���)_O�ꬵ�5�s5��K�)���A�,�VIPWW�Qxx{���\=������7��_���z��|?v�\?�C�V013�Ǝ
d%"(��\���
s'Sh�kCߚ�[v���=�ҝ>/;�z�S������� �N���O�P/X�S�R*Fjаօ���!�=͠h�HWX�y�:�F1�D7�P�Ji���w8�!�9!�Y�����'��Z�	���<�B9��됺���XBL�P.�����
�˭H�c�p���X}�ɧgB>�32��p�R�t!b�1�[Fm��4_�F��d�4�� ��Ԉ��x�d��/	jM�Pm�jc�\�n���&�����ܻ/���O
�z��B+���P��R�'3\�%�[���oFHG&|[��ך�Pwtw&�G�0ra7��v�q}��	�}�L�l`k	�H3h��A˓~ϮZ�`��1BհIK�6�c��M�*�	2���4�$�Y�fY�(Ŧ-��)�@]�a�, ����l�g��@��!�l�`�y�F�~�!@J�#Ò����=���� ���?i� -��9y2���'����D����K�3�9т�c��Xh�1���oX2;����ϮSCT�B}�\vc�63@�o9F�$���r��O����m 9ݭвЄ.�^��Q�ހ�~�N{J��PR]���n��t;>�L�g[G'�ZZ��׏��qZ׍��Z��d�Z��?���� ������
ӳ���\�ƛWH�&7���(,�ElL�c���3O�7�D^v���_\X���R�7������H�KA}}��+��Ĥd����N���p�"����㻿~�o�����s��i��X���6������k�rqs/��N�t2>�<���m����X=z
�n� -ih�OT�=`�l^JU[	�2tۢ�[���N�΀�MV�p�=�F�i{0t�,�wB	���D��n �>Ҏ�#m���@� �PΎ6��\w�5�Q�J���0t�w��C�]�D�B����ڗ�l�M�T@kP����u����oF3����0f���@;мB���y;@'���C����ӏ�D�$Up	�<e�r�t�
�о�c"=��93rW�N�#�rgD��P΀>�����Kx䵇q�QI'D��r���\��g��+�����\WRW���+��ކ��z;B�Z��΋�������98��O�_ ���"������ſ��{�6��[�F�ui=���R��*�t�������;����G�N�6*�wѹv���*��Y�o���Up��ϸ�Pp�����(�������#|���iݝ��w ���'���I ���lT��c3$��d'�p4ɞ0�H)Et�3b�	������& �,��!�^9>�b�.�����?O��Ȭ�@0�����oK�_{
|)������$�ƎW±2v%p���kY,*�[q��Sx�Շ�����K����]�Bb�#2�CS\��,��l �
#u4k��ME�*[ѪF�-�.#L:a���eG�D�'&�5ѭ�Y�s�P	;L5p����Lq���m�p��y�y�Py��>�lp��y����,q��y��hJ�<G@���ӶX2��a3=�4����%�匮"f	����pF�h+�ˍ8�)suL��`�H	{���WK�շ⠮)jU�b��F�uh�T�ުt|������{<��s%خ0��xk({C��Z��7ǁp���F���j ��0]�bkޟ��Dh6���3��L��6�������1�}Lhـ3����l	#��B�.Z��ϦH�r�HXTE!c���S8r�>��=��<v� Ν>�C{�`nr#�謯BCi>*��i	(H�FN\R"�0_W<<��nOWkxy����N 4)9D 4=)B�	QA:[	�CXٷ�������g����˟��<x� �$��y� (��6���ϕ���BMMIT���X��:,�Kd	6fܛ*'bK3I�\�'����(����Hl�eF)c�3��PΆ��Z�����q�PiSFc�����?!C��e�sc2��Q^��h���QC��c`2B������6~-#�;4����B�3���Z������-�r&�3��k0��qSE5]�<2��o�25���� )��긆�z���C��-g����Z�2㒯	g;��q���z
HR��ܮ�����()�5���z�>|L���eޟ�'�t�F&F"���|
��@yjfa*� uvu��A��7o@aI~�o�����}�&n<~?.^9�c��av�(��Y�	��·;��[ �Ё i�	=+���� �eK ����܂���s�
nLr$ݻ#���p_^��U�n�'2�[�5��V2�:�s5�����L`��ଁ�.�⩋-���衍��Z��]�\԰�A�z�b=��*Ǘֻn�:7y��U�O�ձ�S�di��{���:4O�]���]U�_祁u�t\~=�w���
t�wS�ut{�z��߃u��Ιއ��@�9K��x��´/jt/Ro�z���P5߂�>}	O��3����3{��N�74�y�P�4'����0�K 4�%����W0=��1Z�}?=����E��Ndϔ �%��^0O�#��w'�
z���%�j{�B5�FU�U�Aq��&����Y����w�A���W U�g���%c�@�<�ܕ%�F@fJ	�NT�O�(�R
�,�~<elJ1�o��J��cL@ӑ0���]%�.t@�n��[w��'[PM�=�":�cR�J��Ne�V�%��{ύ�r}�	*�QM���?���L(m=5�&��un-�ݜe��[��F�s+�-�������XXݍ�=˘޾�p7���9�:�PQU#���|WO�@hw/�5��J�z��ki/�
-���904�}VGEF�U���b�fy��HOFJRV�w���4����Q�65)�w��Ϟy�c����CMu=rr���H�)���9D'�AMG�L��K��w�������/q��9,.��������l[XEu=]��~M/�sh�t���k�Q��-�r?ƶ�����N_���P��N��d�������t�S�Ѐ��2d��G�͐Ֆ�m�-���z�7�d[ta��4�/�Q��W��k����Ul�Qu��@��㴑���@���\�\���SX�o	�'�
�8�VGE��z{�@�;\���r�.T�r��Z�jz}��f��k�O���h�X�4	�v-K :�Զ�	����m��_�؁��":|e"��3���З�������N���4!t� :{a�t�ݢ
�G���[���_ƃ/?�����=�yy�Ȁ���
�9?��k����듒N��2�\���w�c�:Hed�p<N���J��@i��g׶�'�)����#�Jy=��t?	^��<�%o�s�v�t^m�/C�C�t��RI��^����uIn�i!�qgC�q[��ci�&�Ru:;��N�==@�['���r��ͧ��>���q'>9����α��g�u�E����C4��ay{;O��c?���6:�N)@E�� ]C�4� ���^��ƕ	����8][���kJ7Iާ�0� -� ��  � �ЙTL�,	Dji��$�x]|E((���PBel�?����G��C<!4����]�Ý���VB(G�7�	��ЈLW�HJ���h2�����'#T 4�ێz �̜��(�_E\��㬖T̮t�̅y\�@���H�
 i��[}������wg��"q�9;[3P�4ǻ#�&��_���>yo>]���r-��L��㔆Y"�L�Z���SA��"*�dQO�Q�A����nŘ�!���\�xXa�P]r��'��)o�6�݊�:��༵�*/�Z���%N:O9X�䌽�<��єÖ�ƒ@��4�k��"��0�In'jnHa �Zᨙ��a��>v�k`ZC���8�猛yI�Y��S����`�)�����i�aQC�̫���o"�3vZ�g��}YԚ(�p-���k�߾�+?ÍP�5��6d�\��l��_���Ùp�ʇEotZ"�E��n��fk4�"��G}�t29x^�@j@�	�F=�b���3:-�У��4�C��@Z�� �UD {�	�{�p��I<��M\!طg����y�t����%���ICqJ��"�����z#��!��p�����\��N�qF���-B��D4!�~WT��J�EyQ�ښ01>�����|�5<��Sx����ߑdA�k������_��3RU�
/w'P΂�ڙ@-E����� ���#�jo�=ú����֢�-g7��QF��!���Ĉ�����4�VٕfE9#��<Dg�gWn�_oo�</s/���3_�P2�R2>9�H�)�7���SiZޏ_/͐�1x[i�[������:�;K��4x�5U�PAFWSR�r�P���M��9��������)W���e3�^������L�i�%�����n�c"i{M���۸j-g5�c�z��30�'b=��4{�C�p�ZƬt8~=�VR��$4q;O=C=��463�}8�m@�<w@� ����NJ�����Up_z�gx�������A��rd�0,�p���ݳ�}	��F��5v0 �p�kE�y���$�.hTb8�R����ĬxD�G����P�Ӂ���\�!�nYClax�2]t C��쩇���D��0�\�	6����:-��K�Щ�M�:R¤+a�C?����>Z`�=��|o�����=��P�`�M!��l������O�u	���X>�66�p�r��<�k�{<5�����������&�����@�<���0�I�A[�yؗg�6�����>�kO?(ڀ�@bݠ���<o�e8C!�VU��ɁkY8|@9�ߜ ��BW���q���3h=҇�ՈH�oC(��`�j�8�A/H�P/]h�iA�^2$n�Ead�2[�?d@7��T� J���yg0:�(�t^~�	]�~�pK�3=OmSܑ5X���V��V"���X(��d82,9sɀ�N��,F�!j�Z���:!��?B*mۧ�6�%Z�T*2����|�Up�,���ZQs�U T��=�"���m������4m#d�����V�;D���ʓ�T��6��ScH�H���.��4L��H����ltucxfN�����.�o`��t~ݽ�.W��olY��'g?��gk{�X��ك���C�<.2�<K��g@�mhjDUmJ	�e\��(]�m�馲cK�**C���1��W�� �y�}�O`߾C"{��"�� �M�\Sks��f������>.���ԅs�{�0N_�"z�]\>���}�9W4�k{QRӂ��d���#.=��1����F�����!W�9D �$��6�� � >�!��p�����>���J�U9lT؈MaL����*4�jC�B=A�U��@��~4�g�	"R��i����j���9VjA�!�0@i��'Y���#n��d@�V�Q��N�]��Lv|�����J�ɥԬe@Sz���r�d{5�wq��ΫNT�m���l�OЃ�eh���;��I��v	@'�Up�"iP�'Ct�@�qPQ�� (����&1z��H �9;�Y��"�2]�kK�.�荇��ׯ��o?v^�) ��� �ҍ�%͋^p� t�>�QRW��$�RH���\ �I�M9����S�6�h�9y��}���u�:X~���B
�;����ZOt�eFU������'@1�{�|��.����:~���^%hя�������:��@��W��z�����"�L�X��#���A����/�$D��4�:ðD����m8y�Zn��A����"�ۭ�����ۂ���q���L��D��@i����[��/?gl�}�4�,��V�M�~-'�:Д1��:�G�E��*�#��@y��gC�\��`� h�h��U�/2�����g!3���aa�:��Lˉ!H�m��x�j<�2�� J�����DK�cp2@�	�<�S�����'4>�	a�._�Ȃf>�<����T'D%; <�a��hT2wV�(��t
:���h(|i�_$2����p��{�F����U7��8��*.����I�H�/�w'�w�#c��n=�h�@t}��ƛ<C7�/�����g��8]��\��*#$R����Oy�k� ��Y���uE��ȡX]�ڲ�6VB�-!�@r<����خ�H��Ü��)m�6zh/*�`�*NGgMq�n��	��	�glp���)xjO�kq~-D;P�iPI��4q��y��y� z���tp�� G�q��wk�aAC�8�l���8�%OKls�Ŵ�2���b�0=��[��T�M�⬝6�9��@U^�x��*���;������+71yt&1nXg��U�0h�u$��m` �@��1 ��7�A�5j�Po���$Pj,�y��P�4C���y=���1AТm:�OmFmc�|޶!5�C;����{DO���:��n�<���Mb� �U[�Zzؖ>s�C�C�L�F��'�]�� 'k�:Z����Nps4���%a������A|\ �b�����t4�cfz{�x/��S��|�>��|�����7������x���ՠ�� 7G:�=�D�OƧ��L�����VP��M�/{[{�?���:���F�S�Rπ CX52YOQE׀$i*ɒ�yۀr����2�	�"80HT���<�	Óa�Î�� ?��dDJωϑ��J��h����-/�>�u����a�2R9K�YP^��⸽z/�cU�
.Pmu5Iм��Om�>��3��=3�K	6	�4�e�J2��
�2���*��(�l��Zi;X�-��-��o"Hr[Y�)��=�2R��"�����8�:�_rlnSk!P�U���\^6��f��k��v��*�*��-�;'���媸ήNX��^$$ǋ6��N��x�e<��x���^К�b*lƈ6���tΞ�wxۊ(������B Ԏ{��w�D��=;�i1���v��1p�􆺝��W�� [=��Ɛ�5���)����`����L�)d� Dl���D��[B6�
[�^���AT3(�XB9��6����YA!�[#m)l c��D�`K�5��B>�A��x{��%��",�)܂ރ��r�V�eyz�b�-���t���Nl���1#�jc=!Ԩ:^S�p/�aU��5�{
q����^��/>��}��Hð�g�A����N�I��f&}JBn4�-Ud@}�ښ�̱�~�
��=�GQ�T���tu����Vَ0O��~�1�Ì��� ��A�MGtB�m@��>e�C�Py�
��fl�و[6a�fZw'>)8�����u�1�,=�4	]6t��{V�Ȁ揕�mo7*�עh�seb|O�#�S
KiF�h[)J�W�t�R�h�V]���R���+�-�e^�Hͻ���]�h&�v_�2&A��=�֬e?9<	�5GLG[Q�]Rf;F`=҃�h<�IeQΊQy��mT��O�?؎Z*g�Q�q� �K��*Ohy�b��F��'�y����4v�_���Xؽ�	Qyy5r�PY]#�����.B)gA�](����Ѕ��s�
��so����M˚�:l%�*�P^YFǫ@vV���=K���@'!���+�hkG�_ �+j�ŧ_�n<r�u�"�:=;���l��� �� 3;KD%����aay	}=��Ď�=8q�@�����Ut�N���y��H�)�Wp"�SR���q��u�L����Ӌرz��\�s��F��ψ@�z�����zt�PQ!�ʊ�~6kn���1
�KP��, �v�,A^j;7L��B$CR��z��dt�hF�A���T��< ��i����:5J~�% :xh�{�Q��U��P8)h���d�e;�P�D �j�+�_����~��<}�v7�h�R3F�ucd�Z���C3��O����(F/Ma�<������|�x?�^YŎ��qq�?��޼��ǖ1|~T��~���. �̧$$�=�pJ�Ǌ�H�#������&�|<���{��i����P�(���!��<��H�<$0�p����%��4Z[h~��]�Xzf�~v '_?�?���^¹�.�ě�q���8��1|���݋ه��ح��5�����va������~lh�<P��a�n��u��3�M�\��(�M���%qw|� ���5�=DO�k��L�KZ�t��}+z'@oe:���,2/���`��(�	��ex2�%�P���~o�^p�<K|y� hrI��|�Q0Fi9��_����A�i�3�	���Fa1"�]d6�hjy(�K	��OB�]�煈w§+B2�J� �tYPF��4M#��:"��숈'D��"6�Q�JwC=���9�[F�� d4%cr���[�����®fQ��9�y�p��wW�{R�ٝזx8s�P�kJ1�{K1z`o}�~��7�ۯ_�/�õ�t}�c���x}�ś#�r+�46!]K	Y*
�WWB����d�����2hq����9���`��&�6af�F� �.��cII;�`YQ���Gi+�j��j���v�8���Ύ���$���SK��7UwOۘ�gCyJ=������p�@�uq�
��t���w��*��T0o��EG#�t5Ţ�>�t0k��qYLn%H�㨵*�l�iB�uSt0@���^�����~���?�_���]㈭ˆS~$t���K7k�lȠ6�U��P��A�6 
u��P$D*6A����"�ɡRe
�r�XV���� �h	�vKt�C�Oh�k��^�ou0[�P�2���X9�7�|\��+N��cX�N���Ԕ�>'��Q��Cf���j�'9X�Ϟ�ic7[#8��wSC����?��AHO�D&���QS^���:��Na���8y�4}�&���#|��/���׿�������*4�T	���vc��������Vp�p U��TQQ^���H��v�p�����=}�D0􅓽L	���'ST��ԻU=W�NTR����z����D��<1���pV��dAp�m�Qiϴ�Cƥ�Ҭ&g.��F�0-Li����Ǔ�A���)o����wy��ǽ�jk�uD����YOB��	�/A���r�P>g�������J.�S:�=�2��E	BH�|=���A�׈��ׇ�qf���u��%��,�,�5��p���"���׉qC�5�t>gC�"���ց�mI�ka
MM����L�M���)��X�N�{	������ �淿�G���w?|����?tK����Y�t���|�{X���Jd@��*��0�7��pp�w�7��.�����P��<�ʎ�Pr5��a���9�[B,(,������)C����l�5dB-��B��,�%��	�	����!v"�����P��� �*Ź<i9�	�q��g�-�M�G�&:B��E�=6,7,7B����&ޟ��Kv!+�$Ƣ���t�Q��d�{��1����oO�uC4h���"\�	���{x��g����0{�fzC-��V/�2і�	1�KiB:2ܕ� �~ے���,$����&�[@�~T�4!q*��	�{�}��2`g�(�����4�����#��*c�a� �e˽����T�\����J� u��G�p1��P6WM�,m@���HF�Bh!�sN2���ђ��c�[�ZC��\6R�3����ʖ�:��KT�#�6��P�	���p�>�z��� �2b��n�Đ+]�%��Sy���"�VhE����8��È#�jz�a���Xi#����m��wt�~����ض���ư�CG�{����7���	Q�3�]���1,�Yőc�q��i,-�``p���XܹL������啌�r�>�nMKK
�����zT����`{��EtwR����t��Q�$<��6���S����ց��*��X@cG"��Dϡ��dT5ף�������6l_^Ů��1��3;�bp|��ڏ"BhU��v`tvZ{��7>���mb}��4fw��ʑ�x���K�cr�"�����/gZ�CK��u��(��D�.m��9}��8�^�2�0�E��	4��l�ܫ�4��븽'W��Q\*��v��� Z�ڄ��#�pR���$�ұ�[Q8Q��<�棘��wh�hKڴ�m��.��r'D�-���C���<T���I���so��4?qe�g1un�	P��ʳ��ry�����%z�.�uYT�>�7��~���(a���P1e<"�=�#���Sl��n��m�Zޗ`%�)p�x����8�E �y�zJ�z���M�CfXq������2�~G�8��\ƕ���+'���
��c��q�!Bwe���>�rO�ͦ/��Q�	Fxm2���>�ư���������U�~b��õi\��F���$�n%Y��O�۫�JCdS�[0@%mQ�:�v��Q��� *� �\(][�fwh;�V�{}�����l(Ϸ�@�����:!�'��_T�MUpF��]�X��P�P_Ȉ䎄��퉘lDB��E�H+�V��@��	���r%|� ����Ff�	�Fe���kc�r�J�p�OsAL:��{��`��д8>e!p���[�'��s��� N��Ņ��w�ս�*�S�7�#�ٕH�L ui��cM��`�쁐�(�>�_�	~����݇��C�11�M7rs��"5�q�ހ,}U��ҕ呩��խHS݂lMYԘ�a��S���WĀ�:L�݋�[7a��,v+�b=�(V�ƺ$��2����������I*\�&�r�q��Y��y*H^pw�#�q���	�Μ1��;s���֦8͙P#�0��q��ƺ8D =���#�ѣ�7�銞:v�B�U�`����zX���n{]̛�aBo+���q�Y�]�8Fr8b(��z�o��A7<<ъ�~� >y�y*�������������$R�k�ז�/�xB�.���P�	 ���U"�24�	�j�II�A��UQh�F��
�S�0��J�¡�ݶ0跅ð=�Q0����a����jTO��{��Ο��c�e'V�a�����h/-@}vJc#���Tz�F<��-`moKCxZ�ł�i����:�-�`C��?�)�a��M@NF,E<!45��];p��q��r	?{�|F ����?���7��%X�������f0�ώ�aqr�m@�U����3ƚlf�"
�F ���;,8��HW'WOb��urO��ʪ�\�l�׫)��̧���h��xc�b�8r\喱eC�s!`169ʙ@�ʘ�9�����`,J�NƢ���fCy�Q�M���_555�k��XNi�2��!!��xJ{�嶟<��~�Z�y�����700�O�9O��I!�=��%t� �^'�Hׅ�-��H(_+��q)������_��䶞�Q�餿���T~-�����0�uΎb,P+�n���Ն,T��%<6(�?���A"���⻿�A �����0�+��O���k���Oq��Q*X������ :G7��3a��P�����v�5��0,.A����E ������a	��[�|���%z��r�"S���)nEa-��2a�Q�����rQ���u�\��@��PsP�(;ȅ�8�!�A�D.�8\!�-��M�n�s�FB�Ʀ:��:�>�NĽ�{h��p�!��\DlJ���$g�-���9�f.��f
�<_�7�ò ��U���M���{x�g1}�;!
�Z���=�B�U�l7Q�;!����Z����[m@C�Ґ<\���,d��|gZ���
�������"D�6���0K��A8}^P:'C?#(��j�2Ar�zl��������3�n�
+?8�{�5�ޅ!H��C�B���	���Pi���{��!�)'T �^'��+ڋ�+��@�2��P@��_%����<�� �=��Q��@	�Շ�Py�AL�T�z�U:�D�P9�D����>�ң]�?�Y�>ԉ��C���% ��omY�� $.�S������W_��g16����_؉m�v`ye/V����%�N���Ѻ�&��`��w��a��=��	�ph��?�����h}c#*k�	���JT+	�-�1���S�%Y�{���޹��?����%�/���v�!�9w	�I���DAY	r�aO����,mG�@7jZ�@���001�q��Fg��Ge��)t̢�g
m�S�Y����n����>Է��1�m� z ���č�_�Ͻ, �T���`�@��-�C�euTЍ��ᡍ��bt�� ��0A��z�N�����"�I���~Iv�B��d|�T\%���"K�/ :xjۮ�����ys�:Y��޼��[n=�J;!mB�4Kz� ��� :N��+S� ��˽��0,�׶a�����b�ܬ���. }���q��9�^^��0,��'���"<��n�'�&�Pi'D�N�02@9��O�O�r�L� Ui	L��|'>E<E{�3kh���(C�_�h�V�厒��9��_?��\��Ϯ���'���>t�@�p&�	�.�v��2�I�6�ݕ�d��v���$7���A����l����\��?XE�%�����L4.�X>cX&����>�O�b�>���#�7���6��AQ���� m����������
xR���)��n e\r�۹����/�	�m>�w\�(�*�-���-UԓU��Jn��xB��"n��7	��SDh,�@e��:�'w C若�$W���સ\%��~�,hI���{7��� ���pz�Fp>���tI��ؠN�$�FP�rÔ�M�H�@-��K��S�dG�bl� �?uLT�=��-�#�.Z ��ີ���+n�}���$x�%"�5q-�(�*���)<��%��������̩�#*B���H
�C��"������,�cA YY���i~Ju�0�hB�4�����e0��ە�`����Ҕ����{�lƪ��P,S����G	����8� �B���YG\�p�E/�;����ᒷ#ι�����N�>	L'	�ϣF�Fm����V���Ӄ�j�G����e}5�2PŢ�
�),Ա�L��@�0��6cy�Q�3�7Q�Q-,Y�a�^�x`�8~��%���m͸��=�T�*k�UN(�s=�Q��J�f�����\E
%
�l�rf�!��KP��p�Oi�2o�}T�B@���	��0j��aG4�[#a�	��hDtd#�)�5�hn�Awgz:1�׉��:�p�C��(�Cn�?R<]���$ B���0���.��u�d�;§��P�fj0��Up�hFz2S����(z�mm���v-��]��*^}�u�귿����ZR�ǵk�	�0�����C�u$�ZZFl:v��7Ђ�����;!b�q���������z�YO7O�	��@xH8}��DFԚ�3<��E5[5)8-�����p:��<�d�"6:����j�\����Z�_��,�$#j'��ѹH����aV�M�����`������}������w����RpJ�y;@��!}=B##R2��\�`kCX��	�	e`���3�m�T
P;�˙H3�n 7@ȿ�������V�S�	fp���4��>9�)E*]���u�߭���(�{��ѥ��j�:�����e�Z@5�@���!�[10҇���4�DD[鞤��*��<����h'���_�~���x��W����p��*�'�3Њ��BUd � ���p����J���1�mD�[�Pk�'����P,�7�9�5��1�KElZ�-�r[P�P�yYB�A�n��YB��)fY�6K�� � �j9�pFp�WG(�8@6��i���R£"�P1�ʉ.NBf�aӎ�逭C��w���bnNp��aD���H�p2B	��|{l�u[Rܱ9ٍ����N�����������+�ҵa���3�,ɲ%��$ˌb�d1�-ɖe������T*̜N'i�ݝN�:�~�w��S�T��߸}��=���g��{��ך�&-��-���r�.��F�a�˂0��B�y`�_ؕ�³<}{�ҷ����e��v�[
��ʰ��X@@��<��3	��T�v��f����w3
;7�b`v��ߋ=�(�ٌ��
�up�ۗ�����P�\x���{��a��N��
�j��O���&�Z��J�u=U�=ք]��QAߥ �bx�I�z�8PPB�>?Pmi-|j�	�~���-+W ���H����U�z.tJ"-�J����>W�ZI>#�p�׻U��K�/T@*�9�/���z��v5�k�c�PǪ�֍��m�o��_��:��#-7G�p��M��qOI	�)4�$C��ۨ�qy|�&M����MRד�R���v��alb�S;�������@7��E{��vlW1��rl5�k�8o���)�s��}��_��i~��~�s�����>�^������g��7ncuNr
�PX!^k���o~���oc��	��EKw7z�&��?���.l�G�Ոm{	u���I��)��� g�<���<F!��osgo�ʝW0�>�]���w�sdEU����0Ʉ g�͒�H�w��r8&��j`;N����@������p-٥^C��uS T`S2�J+eXF���������(���8:�T�}3��:V��.IB��>@k����Ѹ�J"���M���C��߹F��Q�(s��!��u@?	��h��J	���{����zW t��MB$ z�# }�����M�~t
s�T��^��*��r=7�0@��8H ] С Ֆb�WVO�4
��;n��!��S��?�J"�b8�:6�� T���>�� ���r� ѧE�	4I째�`;��6��I\��M���}���9�>C��f�l���$u\u��z�E0�]K=���2�c�9���al� #X��&�.�p���:N�^K`�Kx.C?k��\?��^�-�[	�:��7�t�T1�M�;PQb �� P��v������( ] ��i��˭��i�>�W�~�Wb4@�d
|r�`^�q���Z U��<��{U��ǣ�\�_�J�*���K�}��QL�Z�'E��J��aɯ� �H����s.�S�'�T�ɩL TR��l�SeT֔E"�4Y�b��"FAfɎt����9�
�IT��$���k���)Vłf-$$Z#�+����������P.KR"�nV)A��I M+�FƦDdzW��A`Q����ܓ�x�;O�ʫgp����v+ M����LCXm&B(Au��l�Ctk>B�RA������ o|�/=���~�&�}�Ns�()b�I�G6�P��r�84	���˰�� �V&�7�G��RT@k�c~�t�A��&l1n�3\>�I{Vo)��-�<'�Ӝ�O��⌑Θ�4��+��x���Vdn�D��'�	1��	���8j�5�W�W���%�J�UoW\�tq�Eg���.9Z㲓���\��B���(NV8�l��.Ƙp5U z�����8h����9K�z[ฟ�Z\Q�����;�o����S�����;�-N��P8�H����J��n���d�Si2��v
,(VQ+���z6e®y�	��Ypj[�9p�DEl��T\��87��[�� Ty5�Epc��&��-C�b44�CwW��1�ہ�6NU��U)ȏ	C~$A2<��!ȍ�*�_�
Dy: ���>���:��p󴀛���,VfD"'/EE���<�voV�11:���O�W���|	���w��{���&xJ�?��?p�p�H��"`&�S��o��S[���͑�i#c�;�!:&���?M�^RoRjK�$.1���H�'H梭��JI;6��W�EE�]_��w�����81wB�76<��a��(��X;���>��"���(	0
j����vvv�2)p)"����D��Uן��OH���D||�T٦q��V��^\xB���@�&�Q��� ;*-�R6��ބ>�ÇЫ�y�R�O��Ry�LPq�W\qÕ2,��MʴH9�G�l��Ը�JR"^��1�0��$�F�Il�@���J�"�v��d�T�ʲ����u����s�g���X��x~��+Yp�|::;:-aam�bAEl��.�pqs���5/�AP�?�k��rsVg�!$��V��~A�	@|Z8Bc|��c*�N�O�@%������P� 7��W�?�	��j�� k	��z���� ��p��Y�,�<����P,�Mq���$��d�lM̳�U���$+��τCc��Y�XN�C���`^J��'�Rts���GX���?,���B�.բ,�`�%<�R�b�ԈFTCa�}���a@��Ϗ��5B��/����P�)�"��(f��)�_ �W�����J\x�ʂ���70{sY���Y�u��k�5��q�*	�eN B��#�M�oK�N��h+��-!�E�%�??�ݧP6����ѕ���To�F��o�@@I|�,�����[�]l�ˍ���Do��.�8'it�>���g��@%S.���
���?3�%qHٙ��t���nTډIM��Պ%TZ��s���j�����O%C��F7c��@ -.E�X*�mW�o>�C��v�"�S\o�5B	��j���ܬ�Ψ�0�@�L,������Q�%�����U{η`�dĥ~�r�u�;��Q�gXs�t�;���#'�q��e��Lbv�$��?����8؃�&����984���.ZS[�j���š��j[_���$���sUcz�(�۬ ��f?����҈��&����:k{�Ut|t?��������@z���U�ȱص�%�Q�m�\hbF�5���ųx��3��|U{��{t���B��$��'Q�އ��[Q��;����{�'.�б����J�fN���;x��<�x������	�B���H�]��8x����vPsc豏-�Y�8'lڅ�m�s�u�w�rw Mwz	��h �|JV7\U������<ר�N���!����@�����1{~Z���}~��;����Z��l�����	��	w�1B��W��@���n��sځދ��I�3J %��Ax��4�Sj�NQdY�R+�������V/��Gt��$�Lb��Fn�<��}B��<�����~��~����o^ƉGs8�����q��)���u̾2���|0��'��{<��GÄK�.���@�F��8�S S R�|
@��/�ǥ?:	�]<�+`I ��ā�-���ևR��r�Zn�!�\+��'�=�?����W�z��m#�T�DK����� F�F�
��C�=�"��i)��N�qBt�G(��(O�F{qt�W'�p��-�>�Gx�s����r�1,�]VA�X�5�Wcs�&����s�.����#��`�|���%�Uq��񾚮�r�aG&����d੽�N+�2h]�lG� ;s;A�<�k�h�Z��D\粲��s��s��K�%p^'l~J�8p6� |�$|��w�k.��q�}N�1?V��-�NW��Y~s��e��;Q֑�,*��{RQ�s%
�����l7���Rb<5�������B�dHk����������a<�6$��2�U+$M�EY/�)ޒ��MI��H����Ґ]�ll�rM�0�P�Ȕ�O�N��~��m��-�X@5����I(޽��+�X����u��ڋ��.ܼv�n�椼{Rx�3]�a�WD��R�ضbD֬E��t�y�,~��ï��7�����81[������t��03�q[�b�e��Z��V��e��-�l�E����:K=�zؠ/�=.�4[�Q�e8j��i#�2_�S�l,KpR_��8����*��۞��I��H�#|ާ<�����<��$��qb'��Nl(�Qn����f�/��x᪇;�R�J��*�������`� WD���Z*9ok�sv˼��y��w����ܭ��dN�D��:l,0��Bn��	ڒ�p��f<�3���|?�����9������c��pz��aWl�$��bE��KݗD�L"�R��`J1�&�֧õ#���p L��dç�����.EeEkBz��W�ȁu�\���u�@(���Hބ�*;�uh����U���j4��FW�~6��޼��I(Dn��:��Gf��}=����N�{B�'H8�[���
a�X�����رg��ZptnWo�S�^���������ǿ���?�?��-���sTUn������O�!��)K�+�C\,6�����>~��@?x�xs/�
D	]��ƕ5==�ׯ��={100��g��έ�8}������Ø;:�/��^y��v�Dfz�d�Flt"	�DZN[b�@�V�C5����2(.�\U�M�M�YJ��y�"#	�+��-�N�@���"..�׻�ɉ������ �}��"�\ �M����M����������Q{�{`e=�B����JJ��1����L
PJmNq��,���VJ�����G��J���sh]k�����χ�x�m��rN9�<O�^��ĕW�V�[�A[�F�]�ׇ����/������d$D&��0�2����6���	l-�`A�0�]��u��Tz�u`b�� k�� oD��ڢ	�ΰ�����5,\�`�a/[%�+��^�|nb�&�'� 63i�� ���IEV�j���Xĸ�<�+}a������`)Apqv�F
%aAЊpgUӂP��Ös��3�a�L�&�!0,%�CW�8���\_�hD_��H���-�q�]�����X&���h,+�²��ƩxQC¤	����~�S�>9��:�8W-�<����#���%E!XR��0��;�b��	?$�,��'W�����z'�Aږ\x�E���zs,,׉�?��xç*+�	�ʐ�T����Vb�r�<Z��W�����S�tl��#�ceJ�Z�U�#tK�
?� �s�^�g�Aзu�b��Xj�&�H}=�Qt�����@��I�3 �~�T5ug�`ja
k�V�X���UHؐ���J��߂��*���nl�Fx���m�-X?�Ui���rx�٥����u� :�W��*�$pV8�ؖn@Q�zKQ�q���qf;r	���EXt����{���v�m��k-��w�E j/���Z{���6�Frg.U�[1F�7u5�/z^������x�r��P:������@XzY�3�ɫp���.����1>E������(��{p��Q��;�C����ǁ~W=�x_-:;zp|�$�A�Z�M{kP[׈��]]�B[w'���`|r]�v�.t8��bϮ=�VE�߼�Ũ!�~僯�����~+S��;�P]W���6Tl܄m�v�r�V�����6�j�v�;�������6Tl���c��qL�ͣ{��4u���#8B�<���S�8���YLC��Oǉ���y�����c��z'.]A�� *�n�ʒl����'<N�0�����1�[��.�W�Zg[�v�ճ�|�}8����$��*�J&�ܽb���Фd7!t?���|#V�Z�O5����[��|���a��jt����#^��i�@[O��~��ʡ��BЭ��@�* �-�(�N�`��:�h�@ϵ��@Zs�su�>݆>�:tÏ�1��F_�C}�0&	�Z�|}��<�2rw÷G0q� �� zS��* =E }��W�ҷ��ܫ�p��,��г�{_��S��"u�b��(���P��>+��G �?�r��]��v��IX�
Tʜ���"�u��:ȶ��6��c���+�Ǹ��+h��Ϯ΀�*g����(`�|��%�@A%�W�
xF��=�Y�K0�kX� @z����f�&l�`�fk7KX�Z(�eY'��-�e7_{x;�/�~QT$�\�j�F0Ya �@S8��!��ن�u�"@Ͻ~��:����x}h�����Oٍ�7	r�'8J��zL/�ڶ��|v�w��T zPj�. �$Aj����c>[���%����O�GJ m�B��+��	���[��đ�Ŵ�mۭ�.ܹ�X�U�����l��lx$�.@b�T	���AOQ���(��F+��!��oL���( `j��������Oκ8�'�@sy����՜���%4\�T���f]�K�r��5Eʎ�Gr �ׯ�����p���=���k8o]����ߗ���+�'��9�k.FB]>�g`��!|��������cjj/�[�Q_��\�X�����˰NO[��`��r�'x�.{CquS!�ý��`�^���%� t�Z,�Q�s��5 ���:|j TW��q��	wp��ȝyL}B�|���K�S��X,���xD�|�[�^�F����+.�������dg��|V�,�y��{��r��G�q���f����N�w�A*�5��R��`�vW;Ը�:�E�v�Z�&*'/��ʽ�x����A��D��G�z{,w��jw4V����aY���M��H-�n%<z�[�m�gg!|�KJȌ�R��r�K�Pz��;�}dr$#�\rO�b��Z�iD>%�x-�g�P}�w������o@���o�ÖME�^��u��P���p�D�H`�����~� (a[ �w�#�E!��n�jG+�@3�$!�p�m,$�V��~'���w�]e}�÷�w��s���ß����(� (������"4 ��H��C���K7O7UzC\/�-�lH+�^*!��Q^�X��U��Z�U�(&K!B_II	���0�ߏ��;���`�{'�M�()*ƚU�ʢ)�$ɅĲ)�b��V�I�x��
x	d�DE����.*�&�R�&%JZ���#��g$Ym�uW\h�BꪠS�ԏ��	���^���pWmp�$i���A 䶰�`$��"&:J���H�P''��@T����Q�����JГ�L���,VLNq����%JaOժ��B�D�Om̦@����وS�[�S���m���
�J���s�̹��}JVc�d���s�5kbD�Z�h��:�̜`f�	 5] PkCX������;��agc
g'kxz8�]�x�8�-��&Oi��|���� '���������
�0���G�!��_�j�f�����t��Br~�	����H�R�.1��#�6���BT�����J$I�$�&2&���,9OXr>wWÜ �ų0Ks���ж�� ZD��y`� �e�\��#�J��"�wQ� c8�E�,͏�y��9F�o�8��EC�ߩ[��HJ�'KyM�8W-#�.��r�����RB2�e�:��ܡh�¶�����׿�&^~�)]�AzU<�}��
@m	�6"	��>A Mi+Gr��KzK1�;7���z�9ֈ�Ǉ�z{��Py|/�G7 ����ܰ	ի��.jk
B������C��!�.�Z� ��� ��J�T�C�O �X�6ư��O�
d"��zFS)�n@i_%�Q`s+�H	��	��$�pAt�ROɒ+���&���b�,�_���}�T �R$��{ː�_���M(�܌�Э�6�=� �B �'A��N��빃�Q}�	���s�m��炁���*9CT�N)O�&����)��2�:���܂]����j�<{s��1w��g��� ��v��ŝ��p�V_C8Y�����6"��t��1�E�6Q�k?���qM�c���(߸c㣘><���}h��CkK�j뱥j+��ݏ��LO�����>)�����1u�(F'ac��66b����Xdf�R��������X�ev�6��&gO( m����9<{���|��O��s�Ch:HN<����U")�r��.�����10���������F��*�g!|e<VPr�r����K�o3��q�z��A4��УI~�ж۽h�>-��H����@��k��C��s��/6+ ��z��:�@�}
@;	��С�S�4��gG�p�K�$!Ҹ�V}.��$��>R�*��jOs�d�ЮS��m�X@@�� _�0!t�u>��B	�����I��Y :r���;#�5��{�8t��ݛ�!��a�gg��y�p��I�7���Gp��N==�[����N�\c$�<S گ�pG�
���P�I��Iᾲ��J���[=h�I%D �$T��Ĺ/����������.@��XE���w),���c�Gx�8"(f'3N�A����x ��a�J�t$,�r��\
]��Уҿܘ˒��LW�"z\�7�~�0�4����� ��F�u1���}l8(Pi$�zD��5�	v!�p���m�"�CQ�^�g�1��&_�A��Q�g�@�v���ᆀ�d����-W2網������� ��A>eH���౪�T�e�*�k�88~Z�J+ʁ�h���b@�$�҃a�[|J�� ���XA@�݁��|�զ!_�@�%a�8�mZ��M�G��ͩʅVe��hˮ�� MP�Y�h�r��� �P��x�
2�Y��I� h�0��9�y �ZBh&'�U�س*�"���B)t�Mˏ���<}qp� ��}o~�&�tGODeS1���"zW:"��Bx5�,D�@��3���p卋�����1��޴��g���@���2@��>j�|u�p�>+CT,�F��f[#���{m�	�F5!��Z���Q��-�t������r§��T �o�xh2��y���r+�W�]���T�oQA��7=\qǛ����
�䢝�����r����Ҍ�i�u6�@�dk�+��P�����{A��Z☍	�-p����)?g�Sٜ�F=?��Vko�Fw[��4Ee�Bu�讃�l?doN�ޮmx������l�_*B6���ӆ�iW�
;�M�Z�n�
K�ԥ�is N�y߄�qN�c���(�GM&s�Y���xlO�ce,\����>�3.���;�{(��!ne�.��q<"+�U���(��&"�Jsi^�W'a}Z<���Q@��h��'b�!P��I
뻘���>!���U !�����1��
vN�p�Ep���Բu���ޅ�.N�C}ı#Ӹp�vl�
3Cc��`���ru%p������(}RvCZ)����`�)�)�XA�]U T;��R)i"P���Qbv�$�k���z�(I����Ob�WQ�����O�*�@��R4@��:�
*��\b���#��]]��xqY T��eT�4�}�G,��^j_?����=\e9*2\���W_Iz�͚�}6"Zw`�dmY�z(뤬��X ?�އ�X/Ś)�(�▫�r�FM,��,kbA%�SkɔVΡb?�	y|�"*Y�@(�����</����Mݳ���������i 5#�ZZ��L���r;8�������\vw��s��	��~��Og�@]�	� *�O7?�6A��O��"".qi1H�NFJ�J$�"2'Q)+H�gF����	w�s��q��Ӹ���	�	י�ì��W
��>*vSb8%�1��Bj�u!c��Z�#@I��zܮ�'PK0x]=9E%1ⱋ	�:�����:�Y���B��WH��8r�1`kP���0��c�1����lJ������Ô�X�&��<%��ˍ�]V$�c����[�Z���
���w�ڇo���㜏+T�q��a�9�nkl7F^%��;���"Ij�6+ �hw%��7�rlA���;����Fh��V�nDvo9���R���}����1����^W����.�dhjcc#¦��5���[�+��<������j,Di�&�nFI�FBd%���J7(7L��%T��$)�R��i��ճo�B���C����!��?P������v�3[P���PLџĢ��t=?�j � *P	���
>/X.�h������ZU�ˑ�&�!�+�Uܘ�Q�����w�N�La`d��ֆ6h<��0�F�����$��5a׎�سk�Z'�y����}j�x�1\�u3Ǐa}U%�
P]��=�Û��ڢ)�Bii;��z���a�~�S��O�����ï`d|g.\T`\SO(jjBvn�36oFW_?._��׿�E���~�̉Ӹ��9N_����a�olGMs'�/����O�V7u���;k����{x���3:����=ss�/���O��W���ǰ�zR��(�gH �ۘR?�����儠�l/z.���r/F_���k��{y�����p�
��P�O�p�z@A��P���X?���; �5���G	���wi]���t�G�b�:V��N���@���%t^c�?�H ����-8x�:#��1J� z>����1��$oN ���~�>�����a§�K�ҁ[C�;��S�s�5z� ��/��{7q��f�N+��}�_�ŵ��`��1�|�x��,���^±��������@#Һ �8�|�/��q�C)�r�x]|)W�H�k�̂�a`�0+B�3�b\��	-��.��7���	,�̛���.Sbh"."K8�-���b��r�\�D�.�2��T�u�8hr��1F9�J^ʁr1̖��Ď�����=�������D�	��s�="�#��sz�`�c{�(ao�ىϷ)�g#P��p�ɜ��6h;�w���j� (E�[������.{POp�k� �,7\��N�7%���c���� �/T=_��vܕ߱��_��m�W,����P�3�`��PL�@��������j+�`	˧d� xTVMB�����
����u��h��*�9���TV� �mFQ�PϤ�P^*��"a�*,r���o���<{�?��+(͵ak�:d�]�亵��Y���<$��-@Bm>"��cm}1�>��[����{�F��(��GqI0����l����4�/o*C��6,��NkCl�2�pT �Z:��L�b7]���9�ݓ��l�; =�~+ z���,�p��ל�p�Y�y�
�Ew���sT:�::`��gll	�vM{�#���Wly�9��x^�5!��ಝ5�ZF�����Oç����,p���a��A�x�?��]�.��3�>7+���@E�-�����'S�DmHĖ�mx�_���=T�<��=��O�Y	��t8�g��a���aS'%U>�z��k�|0ᇷ"||3<Z�*w;�T�C'�LSt>�:1Љ��2?'�B'��BI���J������X[�e��{I,�Y���u(ژ�u�k�A@4-QA��OY@}����ek73XQ����'�x�)q_� W�6��00]�ź:�Y��E�e�Cz��R� �-���r�@o�R����.����$���>k[k�'�!�aƾ"�~�+��k����$C��aJ"1)U���J9P�KM[MmKq��$�Q�.�,�N,�jblQ��P&`%�Be�&QO�Gq�b%������$���(>+4p)�LJ��yyH�*�P�&�N�H�L_�+�������?���3�5��WD�Y���2,��%��uV%�5j��|��)�C���{Ӹ�
Dj@Q��(��_ V�z,q	��Sy.�Y��m�ʱ�bQ���Ɣj]�e9�|�<7�z ��18(@='''�k& � jnI�0Ӆ9�+;'K�9[����KkcXS�9N������-A�N��/��������,��!�Ct|�c�:������� ����[n4��`�6��!0�
��� U��"/�\(;&k�.��i>0H'x �b	�B�Q� h8�T�0ñ<?�8E�H�1	���V��̷��Y���M]u��L	Sp���ʢ�0,.	�R�-�E�0.��w4��	��0\��Mi0akP��D��'��"6��$s,��(���$?�Ů��pw�y� �:��l��m?���?ŏ)��K8��*��"t}:\��@�a�%6�y0� �oO'|�(I%|�>P���*��l&�Ub�l-�ta��Vl:�����E����.Ej�Z$�_��+Q���M��Z��hw,�Y� ��� FF�� jʾdd�,��k��!�[3��6W%L�8�]hi�F��z�H'!s>5�)mau�(��z���ϲG�,&x��mA_9r{K�C��@Eʧ�t
�6��| ��Nx6c��V9#n�-��)I)�W��t_-!����P�*����K�&|��Bu(?{���#je$���_��c��0>sC�ή^4��v���m��_-���̦�V�q��߳�u�QY�v�ُ��V�%�{�H��,]_��-��ukj���N���S���x�j���!V�����}��������S]�C33�FCK��+��݃�����:NΟ����&p����ƥ�wp��E�Bc{/�5���N/bl�$�t��{T\h-����`r������C�=2��s�q��-�%�>{�}�Bžm
@���8�������U���.�]���8�]���Q�����I�2��Gc�* *^��������)����j]qJ�Z-���?@w��G���WNh\p/�+h��^�*u@+z7.�n�9v�U"T���X:�7�c�:c���F��ad�:��T�����2�� :H���>�ob��8&��w��������7��[�q��1L@�$f��$N??�[_���W��$ ��'b@	�����PY��8/��}���Ѵ���5��o�c�a\�����M���ʛ����!���ׇm�	\�l��� *Rn��$�>M��ahD�$@�������M2��z¨�r>����o��j�r T����l���\�_]=«>S�GOҎF��������(�Qn��� `L@��zW���F�M�p/O��� ��_�I�`%��@��AL�?[E���@U�'E,��o+�s߹&l�ށ���`߅�^9��D2�}�4+UVP��k�*n��������r���OIR$���4�8q�-���O�,w����RJEc�K��.X=D�~��HH,��xPq����y*B	���'�t�@�dʍ��E�4��)n�����K�@��ς`�QI/
W.���b���k�@��$Wf�(��В��8v��ߚ����:҄�7`u�Z��"d_:b��>��T��fN\]�(�TmD˱&l�@6�OnM
��OCj��]�`���"Ǆ�Pxj�M��� ;����=ގ�7C�r�\_���b�=f�'(���`^�g�X?� z����!�� -p���9+c��w����)��Qs���rt/Z�q5�"0�bފ�J`�hC���`k� TA���
�̍1Op�����p?-��s���>S�w� :�`�>gsO�LR(j\̱����V�ʃѺ��;Qھ9�e��c���6ۄ����Y��4e��#d~$�O�mC�Vï�a��`��dq�t2�(Ro�Y+`��[��t7��n�'�Se�Cg%��r��8�K3�}�7,�O�	�+����6�����>��~r
������`d��#��a��'"|\��	���[g;X{Yc���-������� U?�'��^����YY�YY9
쩰��v�|33�g���z��V076�#K[Â����ي�'1�������E���A0!4&&F����X��b%���N�@���$��&�	(
T	4
�Hi��K��J�Wq���dZՂ����d��Kl���fe_��T�'5�)P)`��tJ�#����wɵq=�Z�	h*�(�K T։�3%)i+��͕�� �r��L�,.�RGT�_��7��%.�b�sv$d-�\
PXʲl�Z���و�S����VaM����ܧ�G R��<#Ә�h���*����8�{�*h%|��\��[����
�Y���Cx���s�d��4��ژ�ؚ�a��Z3�Ö�w�5�5�	�Ԕ��2s������t�s��?%@ʮ8Þ����V�Vp�>� �G�#0.H�ڮH	�wf\2�xZf�h�y:�g�@o���OOs�|��A����a���7'�]��8�W����8/���2�.-��bB�Qq��˩>Љu�RIp��6�:���g�-�N1T.��Nʒ�H,+�R�M=�W'�:qX���EY
�+V�0':	+��q$�:a�PJ�t9�;r����\���c�x9��ӉP��0!;;�q����}�૸��mlj݉�u�� :m7��;�`��L�ܮL$���$DʑݱŜ�*z	t��Qw�]�q|υ6l9S� T �x�
�#�����MyH��R��"�RE0t���2;]�����.�|�Q�X�%��W!�&�c;�mz?r3�s
�ʸL�$|n۪\p<+�*x
�J+�*PIF$n�* Z�W���R��s�
��H��~|��@7+�<�P��|6��_Zp��x
�
�
�jstH�\p	��W	4<F,�b�d̕�-�K�ً��<�Fx��}#41�m58q�F�'001���I�����={q��eL>����5W�6�oC:ڻ��էڽ�j��jZ�ūו[lՎm(�(綽��k�>�ھ����0���zw_~O^�|�C<~�9N�?�+wn�ol�mCC��@;:�ӝ�8v�~��_���[��cpt{�8==
��ff��ӏ��Q�1:v
�.\Wu@�:��� vU�bO���_��v��С9��zWﾌ�c�1v�8Ə� �^'�p����ߍ���\��pX�mF�U����Xn����kp��Q�ܞ@��Q��1��!tPn&5�w��)mUF\��@�^§���J^ Q�����{�F�A���@ۙ~��v`�d�����>l��.��n��Ϛ���%�J""�3/�+c~N�|m\�@諓��V t��( %x*�J��a��`�g���1p��B �'Yqc��a��_9��_��s���Rr���~������?Ʊ׎���G ������TmOO)�"�>%	�V>�74 �Y~Q���1�j�S���Ei����h���˭|�;	�3oL�Ʒ�b��#�4T�<*\�p��G����l�T�9����\�%��N*]��O�%������,`�N'�>�L�&T�����)����<�8x�N�����8�q������K�K��%,7Z]�z�K���ǆ����L%R�I�BP^(
8t]���'0�lVŅ֟'�]�\¸��Jr�64]iU��-}C���jD\n���F��F�Ub�|��%Z���ǽ(u"|Q깭��k \6rܒlǚ?NH���Y,��R.�ǁ�F�Q{\��
@��D�%R�	��n�X>�1��u��*��*T��w6'K�\*�Y�����^��*��OV`� sBE���\�Y��YH]S�����
B��nfi4Ҋ�ThɎ���Q�$#'<�@;�_������s��x3����k#r��u�Qukݰ��E���E'����|�qի���Y-� @@��(8��um٨ؙ��@#$���� ;����>�����}i��!vZ���c�. D��,�������I��8e$o	��留Q/?s��*rJ_Z=�'���;"r��,�q���q���F&0����-�	����_�����0��'\vvWVQ9�2ߧ��ly�Wݝp��-��5�X(�'p~R,p�P=O��3�a#�ۛ��J�L������=�F���zk�"Te%�!)?
���"������[�O*X��ca�+65�*�S�Xrٚ���Ju*,�r��Up&|��!nl\��:���&`�R���$���A?G#��З��,)�Ǣ� ,*	 ��ci��r�ie�j�����]��m�p[��xD�' �(qk#����HĆ>=-T��\�N��֋P�eKX����
֒=4��Q�p�"BE�F�wٗʻ�����Ao'_G�{����
f6�0�˦!�%���l,�D
��gI<$jfA�X�����R�8<�=T�@B�X�$	�@�X���(˟@W����Һ�*������� R�S��5���485V>�K� �6�Q,v�Vc!���*0B��tsUkW��p���$"4)�	���BdX(V�$#:*BA��~
��U,��Q��7M�\O�3Q.��yb)��>xR�T`Q�OD�I,�X�X&�n��$�Uܒ4�89��J�7�s�mr.yN"�Uw��j\��U����h�i�+�:��JYe!�3��h��pM����Ywº$!�lc��f6M�Ǧ���``gCG�7ΗN&��g]}�w�kc�FF0w3W�<mV��j��|ٷ�,��jwSX��%��a�
8��Á�\�|��� �$��)p*�!d����j�K�[%�u�T�[s��E���6��|�3��{�����=*MBNs%R���8��)+`[��Mi�<�aY<t׆A'�:n��q6��P,�� ��ô8�IXV����ܢ�9j�S���!�dk�6�R�y�%@'�I0M�Ij�V��mm"�
ґTU��둵c#�m��ӊ���<3�CO���{x��x���ڻ_�[_~_�޷���� �}��x�_�;�x��z	y�+�&��6&�nSl8�Z��6�}co6����X�����|V�[E�w#*�w��� ��	�<ӄmT�7�܇u��	��P~h���s�+@ZCR�Q�ף7�bEJ t�U�x�I�ϵ�.�a�E�Z���&�
>��Ȓc���W��
A<�:u�jv�ǎ��Ve-���^���(��+�$#R��l���|�R�X?e��b�R+ZL�, ljEb@s>	�ٽ�X;X� t��N������� qY��.7b��F�Z+�6��!`)	��Y�S�ڤi��My=�n�׸Li�̸�Wt:IH$z^��V�t��g���Òðn[�N�`��ȡ1��+F�124���Aܺ}�O�C�*�ҧJ�t:���T�ϳ�.bhh5u�ظe;��1�":���m��ڳ���G��}[�m��챣x�k_���Op��]���/�k��.���Kx$z�<�6��1q�� �Oadb���|����s�.)�\IL�v���=�ѩ�*����0zG&ph�$n?z�˷���K�<��Cؼ��-��	4uc��i<x�E�x�
��$Ff��5<�,���}s.����6 :+���p􁥓=,l96�b	��	ǟ��*�<�Eߵ!KՑg3� ��^U�B,��ԕ��J���X:eYłR�ֺ�~$��=���_'�^n����#.�'j0p���.x������ Ov+���V�����=�6�;g	�s�,��ORN�a����S'|JI�ZOi:Ѡ �k�:��G>r�|FyN ] ����;�hYH,�ug}w��G� �7�Q� �胣8F =��E�|�,�>��t��!Lܚ ��#� �CP�υ�O��S�Z���(k���IUV�O��Ǣ��O���h_��zJf1����ů�ǵo\��>4g�3��a�p��Ŋ(gx����Ø�.�l�abA���nD�܀��1�ez�aD����Nn��X�o?O�ZQA�m"���ISc*^&006T�>��*(5�RfAe[��)�F�P)F�@�Rgh$u�4V`%�CvlcK]XqRv�w�O,��T?�BT	�i.j�A���b��!�]�3�ԉW��$i�/PeO�ر��L�X!�|U��y@��o�Vv�����<N �^�@?%��VwY�����R�E�o�ѣ,��/�+ �d�m���7���ߑ�%���q2:�ɂ�v�s��W�G~���h�&[� ���X>B��s>�Փ`�Y�LB�d�]]�U�!l�lf�$��gE�D�g� ��T�s	pfG`�X8�
�J\�O��"��0��V��b�B\����)B4����:���{p��{x��Kx��;8~u{�v��k2	��m�i�A|["���\��}��z�
��y�m�B��|�w��:9y�O]��]�MT�v8��c��� ,n7�C��#&\1�j�Ak�(��Z��y�Hw,�)�W�P-�
��,�(�iN�'�V@�p�R����QN���1�L�,lp><��m�w;�����]�RP��X����W �	������jc�붖�Jм��?^_���㲇NL��p���I(5%�����@(���q��	sQ	�B��)��lPh�瑳
]5����D�C�����mH�3>�m�0���XTK�M�[K.��}Q�C}�[��S�D�>�ՙX���U.X��˸�� �iY�ϖp��  �
��8:��2J��]�ϋK���,&R�t?A��wڝ���n����u���S��X�`*���pq�s�3�p�0�a��C������L�l`�m=3,w3ak
}O3躛`��t�N��������[�Ё ak}3}��氠bgei�k�
B����+�q�$�/��6�Q K ���G�|�)x�@EĵV>�J+�s�4q�a
5V=�L`R@T�J�J,vk��VYl5�_�Ă�19N�M�tJ�N)����R�ӓ@�OR�;��<K�0�?΄��)�Gc�Y�bU�uh�<��)"�b�� ��5i,�u���{��� ��?�ܲ�(@���1�L�>��)�)�d� ��[k��e��C�)�e��/�'�+���)���z���g�/q��oXp�3㼨�����nio���ΜG9or~3���y�L���O�a�cCW�K��r[��=)e��Fд!�Y;�"đ�lc=���x�%�й2�y��HGPE�ca�	��0U�S2���8W>��(��n�4?�2[N�`��8�Z0y�^��+8�h{z�bK;����5P�U{J�.6�Q�*��YY�f�B'�}�2��r��N����nʁQz0��c��$�/��n	�L 4z�b�>�����m�s8��W1��w��&5˂\���O�U�����|_�Տ��[��o���ſ���������PiŴy�5"���?����gx��q��C�r
aY	Xh�88q���$\W��:?Vفٞ��z�]E�R���tUrN��;���w�����n =���F�����[�U��V�!��#���J ��(u1�C>� T��ѧE,���&��[�3"������x$nMG�y����m
@�{�#� Z�S�ҁ�M��Sb?��P�Rm��ܒ^�g�X>K4 �W���P-�J"��
�J����g��VT_mR �w�A�dR;�B�r��|>�� ��͂4p���kZ�O@VU6���Gw"(=N!�����h5f���o�n�@{_��Fp��Uܿ��f�z�SYEG��S�>rǎ��<�s����b׾B�n��Ƒ��[]��6`�����&�vsy�ˊ0<:���{��?P���3��xAY=�^���t���_��;�apt3���?<�'Ϟ+�}�>�N����Y쭩Eu}tu�gx\h��$y���H,��/�ęKwp��S���os�y�YC�o@�����G.���v�z��]<z�9{՝�{n@Lv*�����I���W�pl9���'?�c�6��)�4����ԣ�U��Z���s��)�)p_�]����b�^��:��{���Uh��!̽q�7���at�VЦS=�1Q�,��U�2�[�a� �� ���W|�7}�b����j�.�@O����a�B�� _A�����AB� ����؁�$����w4"�PБ��0� ����Nc����}rReǝ~pSl'����9<��C̾~�F9(��1�� ����B�*p��8pG�i��B�_��o]��\TI�Vn��C�l�p�6������5��`b�Cs���?s3� 1#��41���-<}ݰ"��1!�I�DXt0B}��j���f#s}5��{�G.F#sc,�5*�L��rC]*o�05��g���gLH5"�E� �u�5$H�k�K�u�o�6���� ��Ь�	@ʦdl�D��V?�Kxg�����&�֕v4_���g��-_�뚸r(w��9�5�j�5|)DB%���勢>�WZ�,���2h�f�8P��۔���g'���Rw�I\Mfw*� h���DBe4QY@5 ��ʰ��m�~&�ji4{��,�,�P֮#�KB�� �5e�
B�:X S�|�>�TPZ�Sq�Z)�*�P�Q� ͤ����^���y��H�k�ܒQ3ցW������x��C̜¶�M� 	�� ���И�BD�!�%�l���Y���,�Ol����((GB�)헠�NU��M��Mov���b��~4�S�>�1Ġ�rb=b�����4��N��b�d�:�9 zBo1E\q5 �\p-Lp��l���8bd�a3�	��{{��7GO��/�|���W���u�>~1w?����y��u�13+\���es\�bz���l��fR����68.�l����"�ѳ��3���8�l�㎖'hL_+�ś[����������sG��)�]?�̪\8%����Nd��ɂg�Bf�&ӭ (E@Ԫ&UYEm�S�ޒ��BQ����m��r�d�bI�����_,)��b�"q�)�Vc�\L�\B�\\D�TP�-��YbH�C�2V�S�/nQ�\����X8o��siVP��\ו��Do*�q�E��#�a�e�XN���2?,�6ŒfXLY�g	�@,���hyY�5�X�0�6��
v���%�Y�q�4���)���V�� P�z*Pϐp�S�*QDD��xjLD�Z��,�����i�D�� 5��~
"<�d���
@���*�(5PbZ�@�@�@��|��C��"T	|�H=��P�/��eY���}y�"A��y�[_~!L\s##�O`�|E�U�[2�jK�H�[i�W�\���M���V��4aOk��W@M�oUbE��"r�r_r��r�����K��cey��sj�/�$&T`_����������|�z�F�=b�#U\����)�	��	�H	|Z;���" j��~h���>��Ɋ��#3Ω�0�R�C�Ա]'=,r5��6�.i��X�U��e������px�!jK6���E��BD�ȅ��h��V���*?�ṳ�`�,�!�0]Ö�	*JĖ�=8��<������IL_E�T:��{� �N��;��������X�0�^f��
���iƗ����'�����_�}��q���0�j,�����gy��F`yY��$H�(�hŵo~?!F��y��pJ	�"+t�����{�Q�_����w��?���Ͽÿ��7��?�=������_��?�!����?��Z���5~�w��O�7�揾���{W�^���W04;���8����X��XX��,�AU+�&5b%A.�m����з��vP�mD��4������2h���9X�̶bd4 q��mI��� ����^��ƄP��k u	w$�F 2?
�S�4e�l͓݁�Q�_���r��ʔ˭�f	AY@T`� Tb@U"��������)����m
@����P�����/%�����υ�O�)"����U��EG#�J9=��S��X����^�N���������x����FP���ǹs�����h�������E &��N������;@����މmܧ��'�]�ء��O -((ท���JU����q�ڽ�p��=ģ�����W���7125�=uu�^?{�@z7>Ĺ�WP�Ј��H�۾�!LNM��p��m���0�c[P����~���	ɇ���ܙ�8y�!�����u�p��B�Q�M������y|ϱ#'0v�8�O�Ņ�w���������ނ�-�����0�k.�O�z�С~����8��Y�^���	���|z��:���� ��)���n�b�eeǅF��o�n�y~>Y�.�cG_=���v�U *P��3Մ���@�b�+�)���s�#�P=�m�����?Ё�F��}������ڸُ^hϧ t� :|ﰂ�t��"|�7�I����	�x�$��ey����<�F�����_ ��T_�ѧ�p��1��<�څ�u�p!t�'�aE��#�a�j	#+h���d9�q�[cCS#x8; <�1T���Ѣ�B��P�aT*BV�Ϟ+�U�s*�fv�0����/�R�ܔ�;�2X0�M��X�T����X�UX�e��*.�F<F_��ll�\�2Њ���$52\]�0�׃c�B8YFq��\K�"/��E�؅�W�b��(Z/��p�j�3���fh3_ ���;}���\{����D ����;���F^
)��i��p���Oqk'�M���C��^~�� 豝X�]�b@@%n��$,%�GYp�$9Q�P��j�#�(Eڂ*�kav���JMPJ�0�kp��,VR�
����ǖPi���^J	Q����f�U����V�@�ұ��q�I�{>p�^���<z����;x��#�jF'��*�$��ٔ����*E(�4�o�!��+	�gvb��&��wF��VY-�:[CT�B�Gv�b��1v@w�㠛&<l�o����ʣ�C�8��1� �XA��$���Y@>?i5�]OW\wu�i++L�a����3�����ӗ�O������}�C��_��M��?^}���$(�b�����p�@{��}��g��0O9��<�p�IY`���H�鼹.N��ⴥa�'�-p��Y��b�V��o���x�'�/�]}��������+���ۨ�o�F<V��oS<vf��q�B�(E2��֧��V��H 4���T(�����Z,Z�ݜ��#x�xc	T��#�,YN��XR���:�uT��RA)�ȾVi�6F�ds,̫��Hu۟����	۪�T��*')0Hr�U���T���9?�y����Y��r+�L�Y�7̒�a����g�d/'z�e�Ϝ��SQ���W^4|�F�<�	:VT�l�s����l?@E�\���&)�Q*ѐ���X?6��ZB@�Z PF�iU|�I)'��Q`Q�B"4�K�G��
4�z9�@��\��>NǨM Jf\O���X!������@B���� ���S?q�%|J+I���TdT�/@%(���d��R+���4k�Z�}�u/Z���8 
hk-�r�r�bq�����8���{��3R�F�r�r��������X;�����w�3�g(��rr��W�ӂ���z*.�N��������<<�`*VP�s��V�6���f��\f�������@¦l$lσ_y
�+V«0���:s�x�by��Z�0�ύs�g~4|˓�%	5ń�2��Ɂ_UBw����U�\���H,O���O,O_��|��ڏ���0��~�
��.��k�p���0}�F�1}~�.�c�t��aj������T�ǚp����o�������`�ߵ �%���6��O��.��O�����Ǩ�~�'��%�0[���8�G�p}��P)����f����v�>��g�����_b��e�'rlp1Ʈ�V|�_�����x�'_��?�����g���ｆ��{/�������=��W�/���o��Go=���^�3�����p��]�~x���.޿���U|��O�V�nY�q�5@���!��Ʉ�4��-e(��D�܉̓۱s�����V�@7�ڇ��ݨX Т�*���"��7���X�/��a������ �Tp�E8�_b@�6�"mw�w�ƺ�-�4��# -�&D�T(˧Ă�r1!T��3-��9(	��)\I@�� �S�� �f�m�G =��Hk�}���C� �3�R����'��p)ɇT��������PK0�[0|ʾ���"gG1C\`�c���L��7�=��Λ�A��0��gq��9���-����tt�*��Es[��܍���`dz�<Bv��]�Z��@�	��ض�
##hikD��6<}�u����?�ۿ�w~�#���p��=ܸ��Ocn~�_~��N!���������>ŕ7�E���qe��@k�!�A���B|�!t3'���ݗ���w	���7:���Y�c3�����ԅ=��:���#��Q1�7?�w~�78u�v�5!{c	�פ`ET0l��q�f�]d��8�|G����1<� �����Y͵e����ͧ T,�Z ݵP�Ӳ�J+��o}I\p��L��4* =����A����<G���ݩ�<Ԡʰlڡq����!��[ ���+�X@�g���}��x˂���{�~�FKſ�����f�G *" :�) �xx� z�U����9��a� z�x���p�p��s�>����s�] Ϗ�@��O ��[�8��1\��m{�*:+���d'8E[�9�
V~��t�Cu9!OטB�317���-'O�bebV�$!� J�	���	�͖b_?WDG!<�.��pp4���l���@e+&A��p�s���3�"8���Ȗ��6��Ŀ���H�����&0a'61ק�q��U�aA��^=�2�EXj�=�Ű�6�_�;b��_�W^s��p���4�`�׺��g�& ʎ/�L\a;��7�_�̥Pq�m�Ս�>����-e�XH_�N-|j��y�o���<Q���A�p�.������֤!{'�sG
A�@I �R)�Yp�V.����w3��Y�=%;2PL���ir7D<#����(I���F�"0B���,����)\Y��X=�<��p?v���D( ]U�q�ͫ\���9Hߴ
ީA0t����x�ޥ"���G�׶�6pIuA��$$��#�]���%t���#��1ݥH�,Az[>�[�Q�To�>����� �9Io!p�$�m55�v�.N���=��/Ű�bL��̱��R�� U�'�?@�M��H'�B�$�����r����p�/�n:�_;��<x�߼������o��}��G���M����x�@N�����S����uKcܶ2�H<)��J�Ks�37�%kK�fj�'�D�K���j��3Tf�ٚc��̬�ng��p�j�,��h1F����?�1�?����Q��~�*���uqpޓ�j|�* M�u�J�5d��)N���ڴ^m9�ڕ �5.�Iw��,/,]K�V���>XL U���SD,���e!X�����qQ� �"�E�-�L��m�?�����ݙ�yX�kpm̄w�Z��]���(�mD��6����
�3�e��+S1[�R�!�T����`� �y�p��R��x�K���TxmH�����Aֽ8�E	0�=[/��-�,{sX�e��, %P,��|�/�W��Ā�eSk�$;�R$��P�G�i,���6R"Dc�ԔPk�,%VQ��H�� � �@�f���XP	�\��e��0�6�T�:���z1���B�+@H�v�,@* ��QP�-�� �>��j T��J��@�z#T[T��666
B��u↫���Gy{r/	�q�~��c��I
$𧬓�G�=(��=�T@Q�!<����j�]��Ԋ$8�<7qq���Q�[�������`�Z��\�j,�OK���n.pvv����{;'{e�P'3�9��&����
:m�Ba��Z�8w,w�~�3����D�s��J�e��v-��]W�ئ2xòE~�3�U��e��%�)�U�r����ek����Avߋ0��#nk.��u|��o���K���Q*tgoL��q��:��T.���}�|���Zq��8�<<�����1��al3��傌�8�����{x��7P;�[�VyQ�(O�i!{]<!4��10�|�� j����Cx�����Ͼ�~�=��cZ0,b<�[_��s��w�o����s8�����a��n>���	�o}����÷����s<�$���}�s��A�ĉk�������o��7���,��RB��<�u	
@�9nX��87'�!U\p����V��o����`��~��O�U��ҩ�(߂���R�j-�����)@Xv4���a1�,�y��,���O�ϳ���;!��I\I<�+Ӕ4�.U(�L�ܤ\p��7h�Q��Y�#`) *�W�@�q���(�|]ԫ�~~�j-�eS�$D_T��).��/50(�[I>$ )��"|��P��X RsU#ub���PQ���m�ԍ��9#1+�Zjp�����1u�t�����=Y=��%�
�
x9vg/^���>lڲՍ�x�꫸��˨kjFvvVgdbkeJ��T����pD�Ebc�FU����.���>y���;��?�~����o��o}������.���ۋB�@����p��c.S�Ѫ�;��ե�k�uK�!ɂ;:}���p��S���;8z��&�a��<F�N)��<v^����.�QeX:�&�52��ٓx�������'N��n?2+
��`X��+�	�=]3�[b������K'SM?;��gG�x��43�P�?\[ P�傫��|�'D���/�`� �s���֣V����p��F���)em:I�:ӏ]Ђ��[>@�b��"p�$�J)����D��@;�4@_���<�$D�G��ث�(�P	v=�����{H8$��I�[�8  r�}b��(� {W ��)q�|`���賓8��9}�=����q]QV��ƫ���A)����1���yD�|8�����}8x��y��pӃ���;��EVD'|��@��@Z���M�G`�6�%�~ZT2��ٗ����֏����/h6�7�N��0�����i9�Z�`��J�=I��;G[*E�X�Ih()@zj<|�\���@Q����w���P�F�reb$Ғ"���Nf
D��������f95��vt�������'P��{�k��P?�`�]����@J%P<�(�QRcB��⎢k$V��
B�Bu������R�b�H �+�E~]:�u���c�\7{���/�i:�;t�7�?���v�n4>�D��%���M��&��"xj�#�[�|���V������7�¯�!A�F�����5���M�ܙ��m���M���juo�$*(%��)"����PL-"��qߵ���$k(��y|<
6�"�"�P�Ք5��L���p�)CVI8%k�")�dC�Ԋ�g~Ec�\C ]-��e����}f�$)��E	�^���7�D��"�,O�g�?��4�ޫ���7�ãg��yOl�,ac�5+U��Nt	��ºJʉ,���]�ؘ�$Bwbi�]�f�yֺXO�ln�*��m�Эƺ�̉y'���᠓z�_��"�r2�e_��\������:O��dD�R����L�p��>��N�l��%&�'�e���n}c\K���]�������o���~�[�����3��T�n�1�q'[�u��y��K���������T�K�+V��n��Z�+Yx��ϙ�)�ym�<���%NX�a��$�h>�'���値ŋѻ����o�?��;��/���?����N_;���T�(��ۦX퉇�X?��`]�
��Lx�eï#���������râ5X�G%W$��r}��e�B�u�
"��-�R�����nqE4������E�����\V.�<�@\z�0o�����W�+��]���=��.����v�	��k�+�0�$?��>X���i��X��].dxQQ���?8�D��
�SY���PY�#������p;@�F�6P;��%�TY��9Kk��L(�,khPHB���4�L�^� �"��G,}�M�J#�#��CR.%��'�(�K���j��$�@���l�Ҹ�jb>E>�4ǋ�Rc��/��U�|�*���AA�B���l�>_O��;>*
���D���-7\�J�v%A�7�-��@���M�ƔP���K���N���d��w�I<([�P® �@�����Y`{eJ��}+�@���$e���{�u��)��DM�S��}e�&�W,��\�����Ģl'���V\{5�b�u�.um\�dMn�N�ך�mۅڰ�b�9���6�T��`�d�����زH'�D�cQ��;�� �X,�r�./f�,�zI�K�d���o��o/����d,&x�$�B'��k`Y��p�<>���ā%yÐ�F ���Y���C�lC�d3����s�]G��y�';�;{ S�q��4��Gq� �ޏ��������	��BON�f�{�&^���x��g�m�GN,lK�`�w͐��:��c�?F�n}���&zc�>���o�ÿ�!���71tv��ް��Knlٺ�D�;?��I*]���D$n\��K����}_��w�~�_�-���Y�o,���rOK$��±k��/����=��w��!�7C���Qn�-����d^s4� ���X�4#���е-��ͨ܁��U�5SC�c5�ڱ�b6��Ǻ�{P~t�Ђ��(�Dvw�:˱����s�]'C�,VF#C�%T�>��>@%W�aT�|H(��-����u�~����iH۾+�fcm[)Jx�P$%X(*�-�Rb@�z�)�&$zQT��Qq��&�s�ҁ(���#�V@�	���2������9C/耲~��{/5b�E�z��Q�[q��9ߊ��*u0�Q�v�Y9�`#�s����sqY<�D�+��gi�Ճ�G��w�	��	�N�CpJ(��ڈC'g���'�;;��A��v��@:	�ݽC�<|���D)�8й����~�����s�ݟ��._��ݻ��q){U&��w��!k�*�#(4��h�~I�ܰ��w�"��a��w��}��ƛ���~��={x�K8�مǯ����Q�i�h������]���g19�kR.�Wp��%��|n�e{GO]���y�Ϝ�Ա386�Gϡ��0��wb_c�18)�s�`��,N���/�x��hF�έH-^���d KW;�Q�0�1���"X��EߩA\��U2�=���+3h�ӏګ/ ��6ԐYj�8��W5��(�<נ�E�8PMh�>k�5�����j/��(�@�N����N����(�����`%��oŶC{�}zTʮP\p��k t�S����H,�5suh��W.�G�3�R?��a��(F�O`��9�i��a�Q�)�O&|<���t��u\=��=�9L�����"ٻ<!t��azi3����k'�<�C�y�ۓ�6��p����/��mG0�`��1D�w<�Gף>t>�w�'h��D��.%mw��(ͷp��ԋ���6B�X8oTnv����D�l~AZ�4˂�	԰�uݏq��0���{��>	������L,�k���g�[k�R���vrrW��,[��Crbl,�L�t�3��d;;���s��������I(�Z�g8P��uƪ�+���)i�HNKG\�J�d���]{�UX����&�����ڢ�ضo�vmFJf2Vy���	�0�B�k����U\r��K,�>t}�53����rɘ�D_�kD vEjn<2JS���@VW�����0��0Z����;>	�������"%S�D�Q@,�p�����u��������~�+�ƒ� �/�|K�d��wt'6v��6e{�	��(ڒ�\h�7�@cQL�,�JB���$���V�8	�P��l_�ɼ`}"
�Ŝ4K+SP�)���XK��&�fKl(A4�(k
���#�`��89Ri���ׯ��*�9�\&���s2���� [�6
�ń�2^��hy"*kJ�1ތ]�;�>�����қx���m�
WN�T��\a�G��!��w cz7�91�wH;7 a�ZdW�#';�^&�6_�2K]TYb�rr��bl3X�-z:�m��~n��:����'�2_��&�0k���4 lR����9#��W��$�A�,ߟ�����RR�WX��TJ;�p<23=��%����?}�{��� ��?��~�k����T�m���9��Yk�!!Ԅ�i�+f�biL1����\���+�#ס�(	|�OHO�8�w�$w��S	v�P�'V-_���b��+��w��������/�?����e³b�S	��p����mH���l���"���;��<�:�]�D��\��C�C�X������Xľ���H��,-�"X���κȏ�tAVuJ	��!�P,)���p�;�Z�m�p�c�1�߂k̾��vmo*ܼ���YI%=�
~�#t�	�I�dG*�T쓝�4ř�ꂥ+���9Q\���Vz�"u�z[`�B+��9�� je��M�����#sI�f 3sS��#ue
�	���ʪ'�)N�z
x�h���"!�Z@&l%"-5�l�"�� �!�%�,!T,~SW������@�.&2J��
���Jy�p�gDh���^�P5I�<�AH�	�(.4��)񠲏�2�P�L�'\��:d{���dD+ċ�nooMr$;�&�f�ˬ�0j,�Z8�|vW�e?�G�jʱ�]�K P�R,�@�e�.�G>kݚ�z�=���Y���bE�g"�.�ќ�S]�X�h�����	�r��k���^wg8:����Č�i,�l-`ɹ�J,N�0w�����P�0�K���J��x,�%�FSb�.����	nXF ]J��I dX6���n��ya�*�([�T��eÜ`��s��sC���w6������J��נ{�GN�c��4j��r���V�%����pJ�Dh~��0{��]��ٛ'�����W�bS�N��� �Y�q�;x��w��4��57� 	Ӎ�0ڐ c�[F��9��s��ߜȱ%�k��{����{�����}���'��`�ք��@����i~X����:	��x���$^>�{o���ｍW>x��\E\E.���0އϚ�����8����O��?��7x�ޛظ+L}`��VTH�d8�\%yS�
��u�l*Ū�2��/B6A���
��;Qѷ;�֢���L;.7b�ZT�tvʦw�p�
�#��ݷ�=�y�	��Q���0���b,5�S�J�&F�#��Ii;	K"��k TW�z����$x�2w�V�pO�D�t�ڙ���� �:ͅȓ�+��("T�*�ŝ�@Y����BP¥Vʸ�B,�c[�a|�	�J�VS�[�sW>@)}|Nݹ��/R.�uԇ��X?5��}|Vb��ԢB�$�Ib@�J����T���|���M>ߋU�)�'��u���K8��*�Z�����I4]���^�+}�煒�%=:�{O�Σ8B���B�0�p]�C8t�f�����4�F�70���<c3��������������r�''cMZ�mڄ�۶a��-X��6�Gumz;{��э�^.���E��,����o@N~6�X�':<9�w?�7��Ǒ�04q��d���8|�$�/\��+�q��#\��n>xw^z�K7�c���N���y�Y�_�~'�����[ D@���t�	.^	��X�=���	����=<}�];{5�m�ݴ�����	���+��ajgC=�� &?'������$hm�ӇF��b����RĳP,���o%,�?�آd�Y��t�$:߄���V^�Fw�ע��4]hC׵>~<���G5 J�89@�G�T3�woE��n윪��#��5K9N!|�P�O���n�~§��J-Кc�h"�voF�l�g�談�,V�)LF�
*I�y���x!�:�����\ �7I=D���ԓYy6� t\����1zc���W�_�����wg��0�d�����/h�=�xw�jץ�����q����}��#M�(�<���L���"�@u�	u����@��+Acs-v�܌�Ѹ�pl�,Cy�ZN�ְ2��`S*�N��VNԄWW�6w�/BZl(����ٹ�(�7�
���y���O ̬������� 8���NE+.�1�
CtR,�2R�� ^�-'gS�4igE � jf�{����F�9@Luy_��-z�K���8�ڐ���iȩ+��#�ʾ�/�6��A��,y@���(�K�iy��	 %�v��E�=�z,(��|�����[o���v �8�݅��r�7d�d�X1��J"�M��D@s7Jy��@x��T�\�V��TK+W>	��4�SI@	�Z*���T�4���#VӒp%���(tB��:/�stua$VQ��, ���"w]2�tT�й1������^9��/���ￆ���ĺ� �fi�Љs�in ��s�jz2f�#udb9�'n[���=�W��5~�Xˉ��l9*-�U��m��� w/�6�.��X���ᄯ#���#3���|N� �D?@O�k�k�Oڋ憸��;ޮ8N�g�wr�âb�|jy�*��o �7�O~�G����h)�y�kS��6�+B���XI6]C��	.��~��v}\ ���B�I�$ z�˧�m�̈�6�i�0�f����
���2������_�����Ư�����o~�?�ǟ���ޡ�ـ��9���mQpڗ ǺT��E�@9\��`i�eRA�]��^
@���`y�?4 K�B��0�ٯ��--���E��E�OP�[��R���'גFE=ւ���N�L��:�KW{*Y�N%]�)��D{���	�C�3���(	�X�=*�:T?@�	F|�"��-D!4�صb�"��� hP�����SA&�M�SDb@�Wjb�6e�$�"6:�1������K0�Z��P'���G��d������� ������K�O ���4e]$9�#`M8�$F*ޑ��\T��(^�$"�幽�	v\'m !S,�����GX��D
P�����E� uw�'�U��*�(�&FM,�+�P��G݃Xb-�Re�X+5���)�$.���֚dN7]��j��&��������d���B��#ߥ��Z;��DeY'�O§���0'h�Њ���
ζX�����
F��0s�~��O��E�.
@�&�o�xbq���r�$�cI����\�A [�O��c����	�&�aX���kDo�����*~���ܭ�>ڋ��5��5�V'��I�0Lu�n���}^�������s�8ߺ��<F��f�&{B]�j_N>��W��.^��[蜟�CV���`Y�
��$�nN�1[�-��ߒ�wK�fّ�q�������Ͽ�׾�e_:��T�	�5�д,e	0/��eiL
��� O�3��������7����}O#�<Ʊ�pX'�
���Y��������+��~�7>|�ÝȈ�8�m���-��\� k�.>?�sR}!�9Ge6#���S�lڡ tǌ&��Rv]n���u�:���`��.�NnE�H%�@���GVW2�S�
O3���Q�1�����X�>���R��m�r�M��Ú�RT��@Y4���fl����X7�ń���r�
���S,��Uj���"�g>�3��k�Kye���s��S Zz�RA�d��&�2,�,���:�H�d���Z�ͨ9O}�2u)>מ�۟C��Sh�.��xRO�6¦��VJ�4�\�d9f��^�Ý �V����z���x��09=M���aLϜ�e��<���0�uR����ݽ���BWO/�޸��G��{�.��##5Eh����Q��ι�Y<}�o��n_���g.`jr
Ggf1J�lkk�޽�QX\����|+��PFh���÷~���|cS38�k�]Ӏ��V��Ņ��q��+���U������wp��S��t]��N��E\�q���ܼ���/�ǃ'o�փWq��-��C�����@�wt;�k���}��$�E������,L����v*۷��oc�ٔ�}��p��ңq��( ] O�|J̮ȾK��K-�C�Tr�Y��W�*1�b��l�g��b����+=�~r�w����8Z�����A��5b]�lك���� *�p@�* �y��T�S l��׏`�9??���d��݇v��ABh��������؃C�|<C=J���q��@��w���-}~C�G�>���-��m���Ηi�Ӹ�ݛ�~�6�#�x����f;��pҁ1s#�!ARjC�y� ye"J�
�Ch���$���`kUB=al�g{S�X��� .�6�&��p�v��ڄ(�]_��5������JCņ2D���Y��L������T.��f�3����������O� ��T��B���U鄜\��Z� *mv������L%ۮ�����Q4 *�o"���m�e��pCRa�+3�L˪�E��L=?��#h�ܮ T��@�"O�� �M�����E��,y@:;�v+Wl��eI>�P�~{�����gwaK��נx!rK�R�n	��ϼ��(���͉��$- ZP��D�S�
B�5��m�u��"	�-#�>s	�e
@ז>	���@(%�4yR7� ����)�k �*���(dPI͕DG1�����م���d'����Sx��K��O���W��/=�T�l�a@%g1�*�uͩ�Ȟ؋�M���%�vu�U��t4@��bT����>��P���6�E�67@-'�}��fB��&�1j����QB�'��S� =� ������9�5�K����y=�$��3�qG[���k�E�fS�o�Ý�1���=z�P�HG	+�m�qU Ԝ�X���8o�O�4$�
p~�*@��XbDJ�5x��O��R�P��4�)������0����\W�o^������7��o}?�����ܑ��w��I$|[2�w��{O2��3ԑ��S���j��r�����\����%Rz� ��$K����p�RX��`��� tI9۲� %|�B'�:ټ�*���Бx�1�/��u��²,B�j*��+@)��J UP|.y��$]#��Y/��I�X�e�� *�ida��?��X�\pm�����u����W����b� ���J�Pi%K������"j,�GE<��"Hř��~��x�X�4 %"�%@).���n+�5���곸��67C9�
9a1���()�@ȕxO�������nn*6ԃ �I �%�>�U9��+n��ߏ��j�
��ܔ�p@ŽUyrZ7Yh���`9^D,�r�օV�_��0��Z�c��,�Kq��k�XSyv���Yc?a�uS�)�!�kRϞ"�rny&�j���ޖ���K\p���sN5������P;�z��x@�b\?@�z��x��e���+ٿe�W\���X��,�:)S�"��@T,��⊻�:1�ۺ���]���?ŭ�7�=݅����/��y��*��<��_����.�5��8�	��q�+x��'x��'h�n�I���#cO9N���Kx���p��<8?��a�$K��֕0�fD 5ؚC�mK��`�BX8�'�� �@���wq��U8�&c��*ݘ�u�R`�!�U�✱|u�+�p�����?�����œ��������]	�����.?z��E����s|���_�����_D��HG@Q
"w��}c*l9�9q~�ߒ��밲�ɵXY����
Us���
e=��6��T��tb�Eq+���S��<���F��6B_%pe3
�+Q�]��0�8�c�?�v���+KD*A:i[R��En�:��l%xnA��#��@,`)�)�̼�2�u�d��8��
T?@y�hvW)�	��=%*Tj��OoVn�bW�z��b	�R,��V�#H;a���a�UAh��v���M׽1tJ����[Y;U	B�$ �&��l�"*�'5�Y���h9߃��Y�wDpZ6�nŵG�p��-9>�'Oc��e��;~GgOatl��9���=����>�b��!̟;��l�J�/�G�ʕ���Dya!�֠�P:33��?x��η�������=Ɔ���݇��.����9�*�S�~�����	�s�b`l?�կ�7�;4������`C&g��"��ƽ��ҫ_��7�Ɲ��p���8G0=�6�/�P *eYƦ�ahr'������������Wq��c\����Ǔ����_�:��������ۢ�&������
'X��������H7t���/^���zz� :�5�� >@,����jATD�P�"��^�o�_j����w�{檕�ث�7� ��D?:��qz@hEgՂ���@%T �a�sM�$D��o�(7܉�g>��ݷ��>;�w}�� (A��@���Ä�i��'��S *.�Ы��T.��^;�\p�O�?�_���
x.���V�H�����?��퇨4��1��A�0v^]s�'Ŕʷ��$��`dn�$�������8���T������x�d�D\t��dk[��+{���� �8"���<nki.��BU�Șj��EE#(<!��JXI�L�WP(\}������$FF@	���b��	ݕ����	�IIAHt�4�P�1��P��1'rI`d̉ܐ����k�TŅ��,�c�"�#�rS:Vn�@^S�����C��+���IC��P�& *��p��_���M"�E�����o��vۃ�,u_� �I�$�����n�*B��4�HVPPq������Q(����Mb"�P�����w%�)�*�9��W��qie*ʪRQ�1yVе��T�p��)VP�x
p�g��}@��}
@�$v4
��qX]���H��r����-��*����ɼ�?�7��5��?���#�M��(W��}~�<-Nq�Q�?��"�c#�gc�x?]9�]���4]�r��& �|�4\��˱��qa��`�@=H(�a�4_�	s]�O��8y������P��V�+��`�^]���E�'��Lp���EW{\�t�Qt�/C�b���A�r¡�=�T.�ᦵX5�������..�*���
>� z��X`E�W@�2��,�IJȜ�{�br��9�w�(��y�m1���Nv�\����#x��e|��7���}����������_��M��AQS)V�� �6Qmypە��YTd3\����l-aO�/�
.TdQޢ@薅`y���>	�K�8� ��.*�"q�-���@,%�."t.��nA ���)K�:r�nX��J�,��hD�+ *V�;e��I���`�I%�r�ńR}*��)�X�9.�&bݢHr5���P\/��}� ���Y�ߊ�� �d�}1&T�?��u^�/oO�H�+�3��X=�*VQo�x*�	DA� �(H�8G�rJX���z�N�b��ZŕU�N�	�ʱ�-�p,�͈�`��������R�SZ���::(��rqQ�)VPW�zH��%��I�%��"Ч�l��P����N�ښ��ܮǏ��
(��|I`�Eʡp_�g�?A�U�+�j V,��ՖU����X�V T��»|�@��K��c5�Ü�x��^�K]+��Z��b���T��%VX,�F��'�քO;���֪������7P�Ee�L�XfoMV[��2B��O�X@�й��,��*�eY��aC�s�@S���x��������IB�����,��@\���>2�0�ұδ�N�m����nw������e�,�m�r��q}���'�s�=/������'q��a�o�@PI,,��4��l�L�	{a0��mS�
���.�����W�ҫ���G/��{/b��0�s���=2Z�q��%�������7Ѿ=<�	��0.��2k�[�N��	0�����T��ԁ����w~�5>��7��uL�H�{<�l�,ؾ��q���4$m�n�\+p�՛�����o��5B�꽛��D8�m� 6	��8����W?���{o>��Y�!S���T8�E�6?�	�Im5��܂�5�Hh-D��\�V�-�'�֡q�<,9&9�k0���txf�_����QK ��6U�f�z�lT�o"���읁Ć,�
����@�>	��g j
���+�D\}2��;/	�sUn���(�0��KQ.6E�� -�x�z~ߞ���U�����PQ?sd�K%�f��lkadV�w^NY T�b�T�%�J���PR�S|0�P)@�qy-:.�ŲS]�G�9�b65�b2.�꧄�
 	�
�������cj��ўȮ/@ߎ!9w��v	�	z�к�ؼe6l����J��|�6BY��5�_;��۷a��X�j�ꐛ����Tde�����Eۊ�X�ڂ�rdr�����_�Z���b���XH MLIŒ+зv͜.��F]�Ll߻���ǖ]���݃��0�e	-k�ڍ۱��I�:w��xO���ڞ� J�%9�k��Xh
�����lއ#'/���;��+�k86r�_x�7����y	k�l���V�Ԕ!43C}����)Npt������~%�6{c�ݽX��6�����]�*%���H��<P¤2���*��ǫ�}>UQ���B�|��BBh����E��ft���c����:����qx ���De����B����� ��]���X�������_ک t�(�J�Z)D���,8�_��Ԛ���n����<�R@�c��:���}�"}�;_؋~��7��w���# �J�ڜO����}mg?��{?���S���;�$�;��0��-!̒�I�֜Ω�T��G̖ g�`{G;���GP�"+E�9��"�Ň�����n�0����8��q�����@DLsG�$W�$FcAm
3����i��K'�#6!	�aшK�FI�ħ�!"!~1�KBdB
"S�� ��!�N�&���y�l�O�o�kR����/:3��sg̏�䄚X�P�Kh3B�S�n`�� 4"?�)HhLBeg�O����Z�����gMB>�]�,�_��|��}#�.�R�?*����>U��K|���Pܧ9��]�rN�Y�Bp�V��7Š`V����t��S�Тڨ���T�g T�%R�H@��y�L���$����#d��Y@�B�ʞ�|�y���U����/y����= M -%�VF#�*VuÒ!��MH�K�s�D���5[TXӇ�����߳�l�M��0�4N��������'%ӱJ���E�Ș[�׎bW�B�X ��m��'��ٴyl�������@��V�b�>+��1��vs�!P�6M�f �P��( h�t�8!���F����8IP�1�1k3������cu�ӈ�jE��	��g����0l=G�y|�Y*��<�_�ctD��r��^�G��K���5�U}������EH4��q���7-�╄��l$/n݄�W���w��O?������~��/a�-��f
[�����s�0&Ս`f�1i�a��1�J�����9������"���"�A�',jT��� **�^�@h tE	�rW��c�,������yN���ަ�cL�T�BǤN�� ���Q]Q�MB�.�S/V��/p�����n0��������[�v��J޺�!�0�E�~S�LR6y������&�lKZ�S T�#�M �S�;�=%�V*�z)���[	���.�yj�R S��*	5�q15Q9�hq�@��4�%`% % %P&��
dJ�A~�������Z/Q��B����<�+C�Q��9�/�@E�]rHy<:9���Jq��Nߩ��PQ"Ŵ�'��=WYG��
4
hXkTLM�"�T1	��S��@����G��}��Ⱥ�ZeX S����禁�Ipvr�C�ku��#��QS�V	S0TBp��amg��Qa�gD�?�ܜ�Z�������s����X�D>�S` ����*�SBk�	����+&�n��<U-�*�sM�Q)^�W��6o����2�>�a�����s�wf5���V¤*F%�W����h��w���x��'���=���	�(~��!}a�;���^���?��ű�,�um�*8$j�H�E ��B�ynf�A������������W�`Ju
��KB�)�aTӚXX@�j㡛�TRз��/}����
���OY:c�a�D ��hw��F`�a|�������^C߮6	��U��IlK���cq("Z��H��\���E*4we9*zQ�?����0���a���}hfX�ƽ�Q�sj��Ŭ�-���Mtr�6�GQO-�	��3s`:��)�~��� *E�����* M�����,$/-P *᷅�b� � �V� �|Nm�gը:�����
�Jh�����ܴ�|m�V!���@;��~��?P����'�)�i%}^��4֮�]y���K�,����*�STN��f	�<�� �J�oR�H���8߃����0:���2+�q^�狆esp��\{�69�Ç�a���شy'�c���I%���+Wb`� 6nވ��N�[0����Rd��"/+����GcM5�nڈ͛6`���k�Gqa16l؄}����ٹyJ��)(@���67��𚑟�E˗���+8~�4�q3����Ջ���X�у=����ر��
��s���ӗnh���)0z��]5�9�s-��M�	��q��K*,W�>{o|�1>�_p��),\���fү+�oR$\��U t�#���o�[Ws,ݼ>��՗7��)@�\PՇ���?�8�
�}�F�>e� ����?��Q �\�y'�.���J��
�;��g�\t�����d#V|��ulKv�����F4mY�7���5 ���{���@to�b�V?�B7B7a����`�
�]�����T�Q@%��@{ϮU���w
��� ��&��~-�d�9��l��M�����><���<���������P�5W������|�x�]�%�W���r,Y�q������2�pj\��jU�v���A�CQ>��/�{� ^��}|������oKXN���Fc��2��Sݘ����%�O�g��J�L�c�h��S\��
���!����ب@��A�:���N�9ӹ��(?o��ҩp����0̩(Div�=썔��">9^~t<Bb	����*���!��":%�Y(��GvI5Bb�����$L��D<��"����E"61	�9j�����[�j�rBM	�f֦�B���1L	c-�@���� gN��b������d�GMriU��|��j�(���ɼ�|	�����7��I��1�ªQ�STO1���OQ=%t�I����H�\d�� h��X��F>�TnATr@E�"DZ��#ųdV��ς��r�rF*�f��RQV��"n+�g&aS T��D	U��F�@E�͖u�0Q�F�<��l��RE-Ffy8��Ȇ9�0�;3l�C��a�m�F|*�t,�ы#�������:�n�0q�Ge�+�^��I�1�����0
���t���bvZ����`�%��9F�
@�͍0���\c],%����c���	w[,�b�(�4ɛT�o��I4��QQc5��&��6����X#��8E;)�k	�Üw��w��?jLH�{wBֳ2�I+K�9N�9��u%x
|��亜�ܐPK�%p>k��\n�e�E}�zG��e�S=UPi?�z�(���9��:��^+}l�tE�7�����"��ǽ��������O��'?����[|���z�6l�Dmk���eЉ�u����0��M�A�4��>�<�
�[@+�TL�x:t�l����R�s@SYe(�*���t��UV��SG��J������_>��c
�CO�N	�zy���Ṉe���������:ƤBG�S7yT	M��Oؔ\���D�@E�׏q�q�+�P���c�o��%�>GT �wU�iPQ�@����In�/�Z%T�S�S��2QE������
�
FDh�M�����A� UЋp6���)�# �O5mH��U�)�%���@��~2_�J-'��
�$�R*�J8� 
&�r�>q"��])�aA�^	�%���%T*�0\^G��@	�r�I�*�NL�����8���.J^���@���O����Ө�eR�[�E��u���C�Z��.mԐ�)�d=ه�K�%a�rdُ�+��2��V�C�Թ�z+�  *�'C��x{�
��lC@�Ǐ��$g�l'8(T�N��y�D����\�(��Q�#�i)4�r>�k}	�%h�pj-Uc~+���RlH T�QJ7,�f��F8�b�w|����[#��3�*�J�-G���<f�P+�E�u�0�{kY
�L/���[�������Wo`��L��{��%�:C�>��-���l�r!3r�-�#@F�"D�5Q0�ܦD��N���VD¹2�kW��q�Ǹ���{�u0���l/,��	�10���U]a9�����0�w���s���M�~�ODԜ
'���#`Q��8�Y��x����<���y��nø�)pH��Ĳ8�T���,�x�|0��T��L$--~
�%�u��#�����]�Xv��N��>��&:�Mtzw/�Z��vt\XKx�;���}EU%�̃ JN TBp�a�����8�� &lc4�o�P����!�
@r�ߘ���|��' -�BVG9
��R8��(!�F�����|�@e������MM����檐��T�<{�xe��Q�C����/�O�P���=�*TT��ۃXy�� ځ���%W��.��,��_"�q\*�J�*����R�./9�-B�Q?e�@BvG�STPm��K�vq��X{'���_R��qS�6�%i�xx'�=y��/���cعk�lۅ#G��u�,]�-��X�ކm;�b��]�;Jʋ�S����JTB��r�K_.#���,�=d����>�=�+W���m5v�ڃ��*��g����_R���,������>X:�{���Wp��qB�&t����к������9�r@�oE�����_x�Bo�0O����g.����ABr5�$D�4N������ ?��?��'�`u_j�f!�������k�T8z�7��20ѰFlN$��9��ONa�����h7���[�tq�Th��2��Ԛ6��YS���QN+H��\ч �.X�����c�R@K�/w���z�� �B%$x���(��3�Y�ƍ����ۊ��a�>B�T������h>(y�K�rd�k�o��@;�,��T���G:�y���PQ@�ir@�lT z������*��
��9H �0�^§(�P�����%#Z��&�	|~2��ԇ���q�O)k��I?��>9�3��~�s=0n�	�]���1����@-ct����akg���afn	C#��|PgW$���)��JBZJ4b��J�)�1݃��#�l�����H@��iH�%��JM��c�ȘPd�f!15�A��	�DHD
�3K�8o)��,FfQ5���AüVh�����|P5��i����x,<�x�{z#42�����˃_p l���a�~D�m��5�5�jD�����b�8d��FfS��a��f^و����x��,�)�bO�	����N�J��}����w *��R�C)��P)B��ę�C��ld@K�$��)���	�U Z��B(���!�V�U���q(%�V7��zV:�J�4TU�ͦ�@i��Z_�2. �l��6/T�ь��H���Ҥ[�C�,��Ф�$�2P0?��t\�6��P��Ǯ��O��k���&���.���ZX���y�Z���%��J��I�ψ�HI�q<P`o��:��b�����<���5Vs� �%��3��2;3t;ۡ��,�bam7AR��Jߟ��p&��;r�v� z�D���;�Q�����acB��1N�jBgD��18��<N�OHOr8�媀��cV�8j��X���V�9�U@5�n��<���D��0`9M���8�s?@�>`�k��u�%�n�u��1�v�����eS'bY8�����g7^�q/�}���~�����ן᝷^£����}�ˇ`[&��� gL�3��$��x:�����J�+P>W�j�@���σO�����4�PQ@	���A@���.!T7��'�������nϋ笛��п@㜸�EU�Ջt�I�z�Cׁ���:��q���I���V�P�o��m��8��yB� ��+!��M����C2��K��z��"�dJn�T�
U�pE���[	ÕbDJ%u����*E�҄�jBF&�D��O�m5��&<W
Ie\QH5����F ���V��>%�S T�р���P�	�J�bRw*�R�Q���_B��0�}2�f�RI�ABcE�tg��OZ���Pe(�(�%��9�	$�*�H��� T�L��+�)�l/�H�a9�n	a�������5x.�j���ށ�몎-��@��j�' *C��r�D%vur���%\���e�3T�<���� O uV����z�M>s�~J�6���Dk T7n���x;fT��O#\�9V����T�4���I������d(@�44p4�Ƌ=ƹ{ѻk��q��#���d��`XWEB��ᰑnS��`5	=q���8}�<��vC'w���w]�q��T �⧯��;���!7��4�mx}<,De{f>� 93�3�0�!��J��'+�p��5\~�%�|�U�~^�����}m"̹��k�vNBr��ba����@l�2�w�c<��c\z��N�C�"�M��q6�?'��'�C0p� ���C���w��{O���68�����0�2�oG�o�r/&�� 4;	����y++P�U����h�R@W�9^sis�-��C-�u�F m ݳ��/��ekg }e1rV�!�:U�6��(�&ɿ@�
j�1�-�����}�#|2�]���yY��9?�K�G��!p�� 9��-!�
x
��m���;�[窮XJ	����]p�"D�P����-P!�Z Tƥ*� ��.����@h뉥�Z�
���R§�Ů�z���+���PL���u�G�G��>2� Zw��_A�G��/#Mm-�v�_~�;l:�]{���×p��m�޻��ƁC��s5�j+����2BZyMJ�JPZ\���`d&'�֕+x��7�y�zl۶�\T���+@��X���Rn_���3Q3c*PTYA���[b`�z<z�	�k��1�C���nW��ڏ����`h�nށ�ؼz�RA����1��;���J���/��B(=�]s��x��x���p��)�_�euU�,�G`J܂؆x�z�-��l1ƌ��d������W0ts�����Wy���-P�]� *P)�9���F���&� t>��<U�(�f	�m>�D)��������a�Y��u�ތ�Ck�jn[��5��ꙁ@[0�Ӣ�.8�D)��G ������vj5�i�;�. ��}pm� ��O�*�R���l��r?7�s�_��
xjCo��~`V��pѨi2O��\�
�t]$����:�	�؍m����^���"�*�c`9yL�i���&E��聆�sdko+[;�5������җ���%|�<��L���@~^���E�L���1���x��Z��і�DD�{#5"�����@r�?rSc����p� 1%)��J@`h<¢3DMϫB��e�ۺ���Zچ���y�a-���KԸ�RCc�)Ӽ�:i
B�A�
B��B`�쨪��Zͭ������'a���PCK=X��#(% iu�H&��(C�!�٤��Ԫ�
@�K�P��"�(�Z �h¦�@E�~>���[�'�@�nG[&��{�xy�
�-���@�n�3�V�� � Ն�j+�Jߠ��s�QӔ���d�p=:R	7��*��"D�it�S�K����,{@95T��>E�ȗ^�k4���HaÜ\� *��  ��IDATD�n
��Y)���Y ��8_U��_~���^|r�����!�NlS.��Yp)��Cq(�$D,�S�!,t�,Q�d�Js4��LC}�62P
�!j",6&��7_J �p���F>�	l{��"�**D�;��Ǹ��P������FK�qQ=	�4�_���X�y~J��Xrk#�!Drx����4���z�$��
��j�r���p�\���������p��^�zB�	�����^S0s��Ǝ���s�,^}�����u|���x���x��M���0�J��r�E��s�9�L/dyc�U ��S(F�S����pX�P�O�� ի�8!ToB�V�}�Jw/���|�_�\�PZ6�p�.�Y'��,�� h��
���i���9o@Uȭ@%�R�pi&t�D��'���'����̉�B�(��z+��LksB�d~��F�@S�y��بX���#�/��#����S�S�N`K`S`I M L�)����a�d��C�6�bDj2O�O�o��Q>����J!"�K(U@��<C����J� ?n�*�O��ran��r>+ꢄ�Jȭ*5�jj�	L
�iK��)ʤ\��5j�� T�ߘ�huݲ����G�/�����j+�d�`)n�BlE��c�v�s*
�f��R?�5ǜ�r?�0���|>,�z��'�O�;n�xe�п
��N�T��4a
��zh T�3�F9��O�OU�� *���TO��O����"|f.F^��?x�_���Ƕ#�46q�0./VE!0+
�Ey8�E��{j��ƒ�0�pC���wp��;�����=�	������<���/����^R
h�<����.Vl�,i��i8#��hW�8��H'�^z���_��Wc��#��"���ۊ�Y��vl��1�:����������G�������t%N' ����f����X��>z�~�~���o�}�T8��c2Ե6�ĳ�+ u����U�H 4U*�f�0��Օ�Q���軹	ͧV`��V�$�Π�\�� G��>f!��i��Qة	�UUp�����}���
�����/	����%���R��d�i t~6�f$"bn
������r�v|��@JW,�PZ���z#!� Z�e��\���J�i����b�М�d�>�����S�SrB��@��r�/���zb	��@�oyF	�p�e#R�CS`H���RFaSBp5ʨF%<W@��� ����v����GM�lLN��������4��7������p��0Ξ;��'N�ȱ��y�&�ߺ���D?8%=	5�(./AF}�$���V.�7o��*�݃��������⇟cݦ�=w>�̛�y��8�	MoY��.Ey}2�
�U\�7��מ����غ{7������k7mŎ���}�lܶG"ۺ��h���8r��TBr>;֫.Y��}��o�K ���/���p����v��w0r�z��nN#���gӗ�	���=��7;Z�C�D�9�8x��?<��䨛<�'0D[�{-Up5ݰhTj�9J1�PmUBe\���=.ݰ,�|QFOI(�r�͇Z�`+V����;�0t a@��n+:	��G֩�e�;�`�rTt6���)���B�B�
�	��?�>¡���!]s��������z��¦[q��]�B�!��Ղ���Kk����M�+P�8!�"!���{�`+a���Xk����W�q���w��=�΁��	�Q3:��tV-�M�Y�Z��ř�5t� =7���^�5T�V`�WL��Ȩ��桸(i�Q��L@An2�1�c"��;�!qG���&1aH��� od&G"5%�����I���/.Alb��"	������W`Rs�Ѽ��Ηa��H+*�Ox4�Б��AVi%J��00&�\���P��d8:O���ⓓ�S��e��dO��D�G'P*��#,j���O��T;�r�sr�F8k����nH%�k SBd�����P���8�z��� ���o�L>��]�d\L~k�͟�2��X���ВU�QM �dE62gE��)�3��-��V���ZP�\ }
�l�e��Zޔ���YJ-oHR ZX� 4�"� *J�PQ=E�%T��J��t�B�ˠs���7+�م|��4 ZF 従�_4Z�)�)^�l�C]��������?�������b���J�E�$�����(�/��si�J#`+}�%��3��t ݭQ�d�*K4[�a������	dM�ə�Yc�jg�5�m�am��|'vr�^�|�(��J8�'<�J�gZ��K 5�)M����6C�#J8� �9��Ѹl� z��c��?�g��)<t��"v�6la�2��@�3���0�UL ���.���(�s��v�b3�!>�C�w�x�i�+��'�w�,\>�W<�g��>y�-<�s�6u#=/V�6pH�I���@�
�f4s	�� �>��:σO���cj�1�:fB�*ieA@u�����Pe� �#���1�\� tL�a|�R@u���gA��7V����U]�H�T�S��c����q��~��)�% *]�L ܈*j�T�ժ��2O�rE!�S�U]�xMW�)ň�*����q��P���&'&!>6���
"�$�V�����&�<S��iI
RET�e�\�OQM��M#������FF ���<PRSq�$�12,	11�Pm�!�*��,<,���Ӟj\ R�Zj�;���SJ%\;1Y.�4]�h^9G=��D�Y T�G�Q�H~@����>H���wJ��\�A�!�*׭��E�^���J~��+��*����*��2~<&��b
_'�q�������ct@l�"�@��]�����(��|@	��f+�Be��S�S �</@��	uB`m�^;�����ë�yf?A%6	^��#x���$&a[ê0X�;oV��ѓ�0�/}�&���}���[�|n���3��Y
@��
��{{Qs�aB �~@�
�mS��~e�L��$��N�aE�2�Q�ӊW�~�ǻ��	6@�g�� �f���������K5]h]"L��u�/֞9���������/�y]\�"`����HX�ZҦC?��k���;/�	���^��m��s�}�����T[�wV�0K�����M4��P)����V������{e��A,8ۆY��� �s_3�w�C����6e���z�!o�\d7�`��t��*�R���	��S�S�7�Ǉ�D�l����k�"��6� � �PB� �ʡo)�oˇꕕ֪�W��o<Fe��W�]�� J��k
� hFo!J��*�l�����"NK7,b�F�,��7[N ]���-X�{��0���"�����2����v4����Jq"�
�J>�
��+����l/�O�a�����w wI��  33��Î�p��<y�u<z��Ѓ�	|;wH�r����!!)�E(�,U9�Օ�(.F�ܹh'T�X�3�j��ۭ�e��c�3'/_J����{��0�q/*韕 )'o��;Hpܫ�oۻ��dU;:��CU(n��-�/�m�b�}X�u�J�7l���mJ��e[v��c#�~@/�z�O�䅋x��;�⛟���虓ܼ󗶠��
�y�N�[�7&�N�����,�C�����va��s�=��n�7� �N��2�6R�S�9 �/*���s���>�T�p��iAT�sd����/SݰH܅���*���;�� �Q��uh�׫ t���TN��S�����������`�U'��v��@�c��:�h��~U����`;�����z����z�
�m��Q=�F��y �zjk�pU(�F9�S�(�m�՗{�s�`�F����Jlu^�Ǉ��?:{�A�0��C;�vkK	C�j�t�l�maK����	z�ưq�s�n�_��W?���QVQ��*WBp�rSU��Q �͌�2o8:���Ş���OC|�?�c��� �&�#--�	t4�����bd��70!ɘ�7�P�MC|F)�nߋ+/>��=��ց��l���c�_"���阌D&gh 4(n�=��ʆ�N��8O���Af^6��x�~�=!��@`�ν����Fk�=+L����H����%�X��M�j	��0\1���5T���S �*��O�l5��KE�=O!ʘI�o�DwЂ:¦@����J��� *��BqeX<3	�s�Q;;s4�6ŵ�4�%J�l>�� Z직�Bd�<P�F�P*�*
� h6��b	�Q �&!���*(�+��9/��1��)�X���w����;x��7���LMdC:��^0O�]N��b�P:Lf�����PD�Aβ�j�1��g|6��9&���g~��	f@��PO�j�6�jgt�3�f� z��1��8M�s>s;t���LB簉�q�#�A�G�k�D�o���S<�����J)5İ�	N��);I�b�v�N�@�Ҵ
���~�kL��#<>!􈙨�4�6�H�B�`+�t�T�@��G��4O��Y!�ش��N���{�������_~�!޺J �A��R����$��7���P}���>Т�� �/6
����J����k�� �6���GH\m"�j;F��0����Fr�-	�J�J�2߈��1Mr���}�F u�XPLM	�ժ�b�0\�ErB�DRW�k@%�sꔩ����J(���JA"Y.���6�T�LL@J�R<*� ��&4�D��P��8Y�
�%��O琠)&�p�9_�Rƃ	���)�C8�\Oo^�tKBQ�CC���� ���F�p�Q�MTD	wTTE	yȓs���&h˹	
$��	�ʺ�����C�%��r�d(!�2.����ꧬ��_�'�V�����,�� �F����my�<	;��#9����T�yf�a;�Q����_��y&Tx=� ������A���{9j2.�)*�T��TR�v���
*���4d* =��*������ۘ��kR#�����ЩQ
��0,
�a�7,'`��W�xK���X� ~�C��q��e���Gx�ٛ8x�<���<?X����j$@�L�~c�Ί�IS"�*�`�N_�s!���c|��_㭟�ݷ���!cyn��<�q&4�I�
�qV �҃���q����O��8��Դ-�e��$9��!���8�ܼ���.���K<����ڵց��N���+�k_��f,R�27S���� 9�5Up+{	�����l|a��mX@�`ƱV�웏��sQ�c!t>*��F��&�nlB喹��{�[*`0�Tu�2��yC���;P���P��Z���O�W
�4�>	Y��5'��R��^�\�c6�Q�*Cq��J�D<%��n��+Uq����PNB����� T*�Jh��*�+�ta��.U�H�t�)���/F���/R�9��<�=8��*T�H;�(�X�wu ��ǥP�M�w��#*UXJ��P	�m?׋U���wq6�؃���\
��@��`i�r?9���}��Cܾ��߼�w?x�@��k�T�mqY>���Մ��r�e#Z6�{�j��Y�#��᳏>P[[�֥��Ķ;QU[���(�bUg'�w?ZW�DnY)*f4���
�[6����غ{�ꊥ� �]=\��{��m&|���G�v�N@w<��� ���篨D{��T���c'q��i�ɶ����'��?'�^��훱py+*gԠ��1�q���k�4�@�Ov�>}%�q�hX9G_:��/�@����~{/v�ߏ����tb�)��
ģy���(>�h2�{���=S}�j�ON�9*]-Q6��̗��mˑQ =�[o��ڳ[�{bNmŪ�=
@�m\���ZUwƦ���h�ݬQA%WTP	���< ���w��&���n���ݰH_�k%���:�^�5�ˏ�Īm��$��@Gmt��� �sHc��O��Q�ҁ��׉~l��wp7?���׷\1��s��0\#h@W>W\$`����X& zN�
V�X�d9Z	3��
Ȭր�G�=Z-����N�Nw]�GϕA\��*�y�k*11j<,�a���� jE�05�Ќ���vlج����ū�����ؾw7z�{�q�Flش%e�������$�$"'7EEy��HAVV
BC}��j�q�� ;�Q�F���;"I��tGbt�PT����8:P~��O%��@*a304��I�a7����X�s/>��ϱg�$��e*�k�'��It��B#��������E�N��do���������xVT���p��S�=aH�4��3h!ݴЁ7!���1g ���Ȩ�@vS���t���{.*�*�R��M�P��:��ϕ�[%�SU�=׎��σ��F�暋]� x���m	�b+	�������25������Ȫ&����>���(i�ф��Ȑ*�a�&D�VGr�h͐`Y��P�&᯼)��Qʆ��!�R��pZ���#�W�\BmN�WF���A:��,Bg�h�m�4�N��}f�I�!�7GN�t�pZu�R"pC!E�2*��Z��h�7$!�9������x?�Yׅ�<��w^Ó���#;0-9��n�MP��� lZ�!�.�]A0<������ ��%�MQf��E�m���v�F�&g��H���[����b�n;l&�23����X��<��[��&�	�)���5	���q�0�Uk�l3�%d�p�Ґf�� ��x'x���S���$�y�6<j'y��ەQS!�����̞�� ��zU��3*�q�%�$tK(�aa]^�@�vsz���ۚa��z'����� ��Gc���v�^��">��|��o����΍kx��:�1t�a��c	�#|��I�#�����
}�G� !!P�Ee�|�4FU0*ŅB�B��I�����6�b܇쫔��c���ꖅ�UAxj�S'����*���y'�j��J� }}
h���b����;P9�v�)�2l�L� ������fk3+K��iL��Jc>�Ɩ�p�}����S'�e��ѩ���w�� �!J�7o//��#2<!��jz���J��@=���.�PS7@��b(��@��6�'Y_J����g�*��jT.�����s��O�Ҭ3]�v�"!�~+nŤګt92m�d���]2�� U�����Ӹ�}�&�S��NJ��f���8[��� ����49���'�)�$��v��$��7�B�,��rO\��*�U2%�V����Q��O� ���Y�j���\�h��ub
�ӎ :��NS�����s%��Z9��� C+�N����3ƊI�Tj�����OQ�P>�	���Je穄P�,3��N���
�MԀ�(�*�6f�R?Ms�`]���[�o��C|���p����rf��*�VR��&�e�0*S�2o�U
�Q���cΖ6���<��e�~��]8���8�Z �6��ƫ?|/}�&F^���%��/
��(�ǔ휅t�B�4n"PΌWy�c��P�߂럽���9^��}�ya�9���MU�8
c�9l�~	�l��f��,�;n��~������c��Z�� 5H�yQ������,v����?�_���x�����vL��S�<�1�:�UѰʞ~,R<�7S��,)E�
BW;��o���A����xO��b!}�&:ε��Q�kʷ7)�$��l���
Hg�]���0���lF��K(!Ԑñ��Ʋ]�vĘm�1��L����!�Q��6��xkL�� ������Gt=���<D�O#@'#��>V_-�;�Q�W���
�T�m x֩�
hA�a�s�,Ԉ
��p��%��JkP�a~O9�ː�#���rBh��C��"�o�Ub�ʋ���;�T��+��?A�8J�|����M͘{hZ%��tK�)�V���G^se m��I8.�/<N�^��ڰ� ��l�����v�GAҪ3=Xrl�ϯÒ}m��K�{�T�5�kc'.^��O��/>~�;_��_���`��y��2QZ]�����-Eai�
r��X�}���������~�?��ϸs��������_ⷿ���?��2̞7��k1@���/;wQf̟�����yld'ϝǺ�[��m5��lCW�ZlضSٶ��q��	�>p;���G4���Ĺ��r��R<O]���G�c�֝8w�:>��g�������+��
��؈%�Ѱ`&��B$�!01�B}���	��p0Sݮx�`��]���	���h��ƻ;���jBnO�R���Sm��NQ6�*P
@J�	MحeZ�S�F	�u���ŘO�T �y	�+��Ɩ|�F6�wx#�����b��v��؊���&��ڴ}��Y�9�9{9�_�Sk�t�kݹm��k�P�ᝍzq�=�F ݎ�/l���[�P.��=| ���U
@W�Z�>l=g{	�}P�T t��>����Kk	��0x�$}���ܑ�F ��:��u�E!��k������XsM��Ft�<�Zh�b��:��4_"�C(/Pa�/��H�{�q�/M���J?�/�c��m���쾵��p�nsW�Ӂ����vt�l,-��maL ���E��9��׿��=�1��Y�9���ù���Ӄ��`�������U�����T��&�� A�>l����N��dw�L�B�o ��cL �
�GI^
s������+����������BE�!4&�C����KWbh��Ϙ���\D�c"�s�_���!����x��5�N��o|�ށ���� 8:�q	( �斕��k�L��5[~��a�������������&��e�diz��b뽝���K��T����� ������{&a���7�NPQP	���h t����>'��A����+R�='� J DnM�k�QP�@Em̢�M �S�̺h�=�5]�F�lf��i6�3�3��6�P��Tx��T:��t�@3G�cQJ �"pf@3	���<d�ʺeP:%��H+�DjE,�S�=?tḷ�1��{���x�?���o����+%�A`GG�8��yA0�p/ڸ�P�5$#^�,K�B�dK�8���T�mM�����qX�x���cu�`����"���Ya+al����I�$<
L
�jr>5�y�&J��֊�r	���0��ɧ��c<�	S}£!���i���h�-&�ʶ߷3|^��N�4�h��"E���,�I�����k� �AZG,���3�zѠ���\��wuI�/f`����A }� ���?ć�k�o���kx���q��QL	��q�3l3��H�,z���1]>:��� e:��N�R9
�Ϛ�#�7�O�vV�i�R������ V���K��GZUJ� J�;C��t�uS�(U}�&ӉOt#��@i�Q��m� 4ё��t�aN��*d�'X`��1C�'�5�lm	�V0!|���7��ۂflm3~�����k*�=�*������b�	���6�U����
8ʸf譖	|	8E��p
|jBFE!ըx��@%��; �}�N%4�xx�v%�`���i��p�1�%��qQ򤢫T���tׄ�J��E��T˕�ܨ�0D���*��+���I1��3�;)�#�'&p�[�O;B���1�ll�2	ϕK-�ʶ2O S�����2Ҽ�2�u�^
0�}��%�G�(�rOD��R���٧l��h2�2��G�v(��J�^�P�ϢrKU����Ü� ��?D%=�������i�f�I�0v�����	P��f�F�%|�E8+� %|�%M�~����Щ��A���LN�LU|(e�QC�KA��U��0_u����u+�ꓫ���=�{��q��a�6�;�%a\m�&��m�em4�JB`� ��8��Ԇӏ���GOp��Xx+�2�1��
�5y�����]<��5y���5��"��M�Y]L�>�5���C�Y�7;	�K�4�9�͸��#�L�}��wq��UD�f�<�����j�.�0^�O� s:��<���>�����?Õw^A	�$��#� ��ɨ �ѓ`��c���Ͼħ?�
o~�.v���?�D�ã��	�%f�{j���2�>�Z�ԥ��]U���zT��D��L��т�[[�{3Zή�\:�[P��&�l���śP��5{���!mA>���	�:0���ZMX������ ���saD3Tf�v��܀덅��ʀ :㝭0�����Q�H��~�/LW&�%���^]����)#LV0Q�N��F�v��Q ����h��zV�h�
�C�(Y[�|gNW	r�KG!�L�+�+#Њ*Z�J�b���	�.#��@[h�'�* �w��N,S��@�/�|zx	�@;�d���II��!��u���%�NM�"�-'���Q����7���A�b���';�sN��lE}���-�����Gx��kx��p��;��DE}9�U�娙Y���;����=�蓏���$l~���?|��'%~��'x�����+QV^�E���h���QY_��-[�������u�^�:w�z��D��uX�i6�܍�;v�y��$l��w��b`�F<>�7�� _~�-<y�_���Wo�ؙ�p�6~����������g|�Ň�wl/�s)f,�s��I*NGhz4�b05�S�&�a������j��k[���!����va��=d��uX���zf�Nm>���� ��V՜M �T�Gוi��@��*(h=�s%���)9�9�B m;�;n�E����
��CX~�-����w��g tw��^@]@�\�\[@]���w	���kT�r��:���	���J��No���)�J��� hۉvt�t�{B���+���㸂Ћ��KCOt��:�]׷�·Wq�ͳ�ue�r��׆�s�sT�S�z
p
x��^>
�+��B�\�����T`�D=��N��0�7��OШ�
@m�`����5��l0� jΏ���!b��q����22
s�<��q�h�9{��Sq��eHIKU	��w�$��">1������v��e��ڊ�+�����	�i���4���"���)�()�ENV&�S���r�9��H�(C��%(olFTj."�2����L���������g&��q�7\���78�#�ɼ�\xDB�����:��qi��Մ��b�Ls��5��J���ClK;:�v;x�OEn}&2g�b�������ߐ\�~���,���=����*����[v����@KV�"�)Y���`��ա�
nQAS`����M�%p���S���(��P`��˵��A����� 4�`�#Fg^��Jߟ��ҹϢ�/К!a��P6l�д�8d�QNoʀ;���Ǐ�A�~�M�~�1n>~A�oV$,�&) U��L�&f9�����+"��S�Q�`�Z6�������sL�`ap.AP�ֈf��f�`��q���v6Ļ�PK,G�G�����>5 *}��R56��Np}N1	�=e�?n<F���#t@����b��h�@�&ݶ�0'���q^���Q�'t�������̰�0�q�:�m����ި�-KZq��>}�]����q��ܼy_}�!�������:ZR�dl�/�	�c�<���th���|��=��>S����S�5Q0+GCn��1�:�ӄ���_3n+ÿ@u	��� �G #�<�p)�TL$|N��ҽ!4fB����G"�'* 5p��~K�La��س����PP~m��) ��=��9>�50( �KJtz+h H8����Nr(�d�Tn�R�V��y�)��2_Bq%�V�U��I@k���$����>�f�!�����	`�Rt(� &!����TM�i
F=��x�2*���(��<ߘ���*�kn#��>�D���¨��8�SQA����6,V�P��:�i�Fه�?Ql�ȾDٔ�&���IɼaOUL��6ʸ�����F5���)��l��t��{h�^��\�r.r�EQ�Pj��Ֆ�bjj��c 5�5��]�n?�	�P;�)�;�	V0����I�M�f�A���O�J��!��>	�c��� ����{,�s�/fҲ����E^��|O�l�	�UHmr�lD�Uñ2����
D��tn^����׎!eNly��l�k�P�k~�ͪ�`W� ��8Xe�8r
��ԣ�x��������vx'|2#	զ��Lǅ'7�Ə?��_ƞ�#Hh.�}~8�+�҅ʬdX�H�����H����#1&� �nn��m������W��K7�<���0-"�}3�! ��8���a,��<������x�����ۏ�E�^��²,��/:���-��o� |���>~��gbL]�Y���5�p�9���(~,R��'#��Xh~{-J�P�Cp�o�����or�����Y���}���Q��e�g*�ۿ -�U�d�d��PS�$��&��4��ħ1�<�N}KceR�h��QB)�c����>��^:�������	.�7�6!M	
>3:+P�}!�6�AnG%
{jQ�S���J�&>K��˪��٨#x
��omBa�o��2���h1*6֨~>@�.wc�B��6���Jf+�nQ�CH�Z�Řt1�c)�M�\AY�sѰ6%'T%R&r	�ë�	���)��W���r/�.�( ]~�K�����:|�lX �4/��nn�6�ƃ��Ϳ��0�",kFYm)*��P3��e(� |�Wa���y�~�͏��s��!ܸu�Ϟ�$�O�At��(.��dn׀�;w��� �ގu[��e�
q���A��x{��-�q��E�z��8��mP@�a�lٵ[i�����7p��#|����G���^z�._Õ�w�����O�į�{��g_�ɛ�qd�0�V��e&
K�Z���s��g�����m��-��� ~��t
��@���z��<��䩥��%��@E�T
��$���)�� ��=N�$��'|�?Ђ����Ý�-��@���C�(�.ڵ�7/AU_���. ]��n��Y���K4
h�u߭�
@׊
J�\ǡ��T9���n�� �P��0�U|8W�!�|�
|>���<сK�� za=�έÎ�[q��K���i켼� ڇA�������F�)S!���*�HR���T��؃-/nǭ�oc�흈���|2?4�ЗԸ10�Caac��%q��5�&�����ώ`ǡ}�*)�W�?bR�������L,_�
���t����M[��J_�u���A^~fϙ���2L�H��U
?Б�DG������"ąE"!"��i�LKCzj:�â�������(�jBqe�wa��6Ť����ѩH&���ƫi�)�p�
&@b�g�3PM;N�����b2��W���x���򙊰�d��&!0"aq	h\Ќ��,��Sd�Fߌ��	���V���)�H(�!���ih6N�{�<��+k	���P J����mg%�@�����UXvb���v�3r�Aȭ#|ֆ"�:9U��PQ@��Z�S�I�T�ɡV�+f#���h�z�:��t����t�Ua"����� ���� h���/Ο��"�g0�!��BZi�h)�	H�����ұˍA�~�|�n_ťo`��m*��u�T�e�A
R9AR�D���н2���7c����R��ge�}4�f�*���o[e������XK��(��'�I%���P-|S���9.�|>x�F�b
B�\BkGGaQ��V��G�d����t.�@�p��v}����I^�����f<_f^�aއa#�6�&���`��kV:;a��3ZCђ��ݫ����E���?�O��/ܾ��gN���3x��:W���U�~�)�������} �-�� ��aP}�^�&\V�xj��	�
|>����P�O�th� ���(a��PBh�d�&H5Q�S�G�%�ƌB(�S�C�D��,j,�&���v�kiB���66������T�u��'���)S0���6�V��'�D5}U��&�#0*���*$����wV��������'*�l�Q%�3PS]vt�JZ�Uy��*��=��)a�>� �+��K���P�!�K�nEU�%�
p�2*��(��]KhP��Ղ���*�E����|�+�.�%�+��U�<c�cP��G�Q�P�O�E�R)w����l#& �UD��P\X����<IɁծ'���}�1��I��̗iYOrS�i�S��T�L�aU)��F���	��}�BS��j1�� ʡ���0s��>����ᓡ�]	Õ�[QA�4������u��O ��I �&���=�N��a6��TM�!	Õ>?E��S��4�˶$���Cx^�vt��K����Nd�.��d?�d¹"n�p�N�mUl�	�e�0�����#�;��{��ѯ�[?��{�0]�M4FHIξz���k<���8I��U��4f�vF:�J"`ݘ��X�H���LXvu���Z�K��w��+����q� �\F��b��ό� �r],��Vi~�vw��g
@/��2J�[`%9��b�������)��/��_����'�A =
�$ާ���&|���X�q�_f�����	�)�^X��ť
@�;�Q�IX���{��I߁�w+ ]x�]R�?@��5G�g)�|�,e�{���!eA:L}����)5S�{XZ���J��hR�hc��-�*�.[�aB��l#�(���5\�:�5����L ��oIk�6��L�g��&�tH�:��Kحt�"ݯTD	�Q	���"ʧF�{���D�jT.g�%���z�;w)t��v���X�j���ګ��i�Y��j�/}�>��n,;�E����@Uh�n��T�|_�c��BM����;��輶������p��;8��r���5����(k,��e8��a˞MXҶ��	���� ;?��,ġ#������'��� z�����*����q��-�]�89��-���GQY9v�ߏ�nڄN�,j���8y�"��:�C�'��y��'x���m�%ڂ�{�c��cj�K7n�E��7��݇/������c��p�/��#x�����/��/�5�ݽL6؎�Ck0�}!��W#�*Q�����g�7&�M�������U�z�^;�}����� �l|�w����A+���"):4
�R@�)dj��<�Uo�G ��ue>�7�P�
���g�н/�����9��G�c�~,ڽs�,Eu�l��� *
����|�bt�_���+��wM��\ǋ݈��6+)]�?B׍§�������z����mh���\�y2=���+0%���T�=��.o��w�������z�f\@���+W���%g�*��� �u��tm>���_����1-~2��T�!}X8��J�Ώ��i����(���3����Q4,����t�T��vn*jj������a�\�|%��"ל�͘�4����\���#?�����O�.P���F +9�A�0�GG!!.��)���Gbb�Jk�дՍ͘�dJ���3(�u B��QB��!S�uZ0�'��a�/�x��4���	�^���$��78a�M�!�� (2S����Fae�-^���T6�.�q����)B#ی����RA'L@���5�uo�>Lh��}��:�) �������<��'5 Z�:)AH�	D^C��	�� ZL�,��V����L��)J���lX6FK�(+Utt����f�JU[Mh�t����hv�'�������M�J����(�@Jqb�ItPr���C5	� ��`��kǮ#���n?������7'
��aK ��<7���t�`��I�H��g��D��r]LQj55��67@��&c=�B�	^U��:*������,����O �0���0[�
|J1�4�p�S;���!tj��3&���p_g	�216P�N����L�9c*������p��H�_�7"�X%�jUR�QQP��N>G�4��'yMGx��b�\��v���橓�`�-�����FOUNo݄w>��~�%>~�]ܹq�ǎ����8vl��a���8Xd�ѡ��1�:M�֦CO�o	��!0���M��C�h���\�/ׂ��T[�� *ݰ<�z� ���W T�� �K �<9�Z�+�F��<r��`2�c��ZH�s�@mlm|�Ѥ?PK>{�t��:�wPa�S��c򔉐.Y`��	����ZM1Q�
G�����)$����k���eS�����b92-अT(%
,�|����P��c��7M��[���iOaT�p�S 4,8H�S��jBo=T�QBE�TE�F��S U�v'�G�*�֡i_mw+���k�L�@MU��?�$�C�,�D���Y
�	,j�O
ie=�lWQT&%�V�kTWm�#)x$�r�eZ�;��d��L��*&���²�f��K~;O�O�']���Z%�Zr@���0��m�L�[c���&�"l
��'bl�D���S��qMO�3n2��)�O�'K����1��ͱ�~��Ӑ�L��?I��J��
�
t�P
��k�w�)���p��)���#\�3����H���q�P������X8��¶ ���T��@�����x���q�7q��U��)�m��Kcp��>��Wx�?��Wn {����ù>�j�`_��Yp���8��!3��p��;x��O�ɯ������0�����XX�K�ɬ( ��I]��6Y����쏿����-n��*j���,����sQ@ySaE�^�o��~��}����Ho��a*�Y TPP�z\v �7�"jAI��*��C��4b�XC����Z,b��,�J�mٶ�(�҈�]�Q�g��W�cf��Or@u``+]���1��5�1R�j��9U��Čơ)��q]~�L49�l;l�Y�~�-l�l��6=�)�S��^��m�P����Y��.)T���J�=�*�S�oE��:[��@iźzTr��
�����"���UE�vh�u�\W���b���j=�FxY�%B U@t�����z�-�ʖa��.X��;xj�m�*a�Z���� ��Z��'���w��w�b�;'p��S��"N�}��-�o��R��פҿ*B՜J4.h@��hj���Y���K�����Msf��{5>��S�����������_ ���O�7�����ʵ�J�Y����e���^}Wo�ƺ�[1�u�����˸r���_zG�;�P๦�}C��9t������Y�=|;��qB���Wq��%���;��?��:����x��'8t� ֬�@��
>3
W����pxF�`j�ƻ;���:�:�Ꭵ;W��k�0p��ys;�}/�kV_ �ta	}�>���6�V �Y��tt�|�?
@�[0� ���j�w.�NnQ9�����`�֥��9���w���ѺwV�_��C����; ��� *��{[0D �
���^ ��ި t%��|`%T �B{��>�^-�JD���s�����Kp�Ӹ��0t	�W O@����s�����.��B��"Db�ЧE�D}F}�{��X$��� K��;ߧ �����kz�����YT,-���8~��?c�0�փ��)�Z����FO}K3L�Ǫ�n�l\���b�ͬ��%��p�r���Ă%K����H:3�|	��я�{�A��#)-�/U�QXV���2�T!>>�^!�L�"�ӣ�M�D�W|���2��A�!�����
4/^�����
*g":� ��)O�CBV94f��N?LM�$�H>��l��4��<��<���!������`�Ť�?4S���u�t���Ȅdt�~�lx���w%���ȏ�=GkX��b�	b��Q���6.D��!��o�q����߃��Ш���=ZxH�i1!��G�S��* ��)B��"D�动�
@e���V`��zTud#�� Z�@�j�Tn	AR�9U�J	��T *
(�S�>eZ�TL��P�Z�i�)�BD
@K�
�_��bN?P�Odd?��H���Z���@�h��E��dq)��D�N��P��8�׾�o}����ݿ	�2Ba��� �ekL�(�y��X���$�#`��\�Pjg�F>��\l1�3K�-Qk��V>8����]��R;��l�	u��FT�O-|�#�>k����z8C�<�}#�#0�����Ӯ��^k�i	�L�ԸZW�zZ������\�s�ϳ��P�k�������{-��Fd .D�bh�f�X���+��~�L�=y_�������#�bcw��>�:y���C\?gX$L�i��h���L)��1��%�Ӱ<L�r����3����G-�jCr�j(�Iu\��w�	����$�WW
>� ���@��*P���iO�g�TU�e��D�����4�N��.�~�kqL��	��a�a5�fn��
��w���Pa��P�~k�P�t%�(����4���$5�$�J�)��@���@�D����S�݈���2�)�/��D%���U��$<7*\��j�L�I�Y�B	�MN	���n]8-�"x>�ɩ����	��NM��
�U�T1"�<�T���܆�6e�S��ET֓y�~�r�k�Sr5=�=�Q��͉j�&W+�@��V�n
l�Γ�"�
D��.�OL���݊T��m$�V`Qr6P %�W@W��C���{��*��C��]���,�Ҫ�r�r�:��K;���FDD��{��S+��:@����Lv���L\��8�3�n���X���386j�]�M�si�8�0H%\
��9��O��@��T��R��ͭ�i΃^�T����[-�9�*v�᪨�@ɩWN��o^�����^�o�Ų-k0)���4[���@�p�>	:A���qBHi�w-C��>�pw�x�W�� �_D������Y�-�����o��O���[�p��T���y<����0ea��Xg��(�:��5����¥w��n?��л���Y��I�=��!|�Èf��P��;�����V����+|��?����+a7c��a" ^��O�Q�;����{��k�����: G�F��p�ä�8L��t,�u��s��i��������\VA��Cњj���c��f�s��:�೙�#�?%�VBp�%�S(�}�(%��nlDҢ�5t,u�oc S)x�ﷄ��Z[)3�0���),����056���X�5��c]�-3��w�����e�vcfӱ�shv-D�&��`=��%�uG)FT���bi��MQD�Ȑ��5�f<-:TF�|@�
�*|j T�}z+ŉ
	��*W T ��F�P	�}�%�t�r|	/U�)�$��P# ���J,nW!��	���v.:�R�K� ��h˱�h�Jߡҥ�@����<���E��M�p};�.lDS�\����7�I%�H+KCfY&�1t})�*
PT�G��C��f��lýw�o���ӿ�	������������O������ϸx��8���^ē7�D�ڵ�{��F��Z,no��}{p��<y�]|���J��I�e)�l�RlڱK��nܶC��2�ݹ� 6n݁[����8{�^�?�������w�◿����=؍%=K1{�<T��#wfbJS��� ��M���D���*j���s[p��l~� z�oņ���A7���#���K.t( m�@��}� z�/T%���@9.��pr�|U�H*�>�� �<�.�����pv�ُ��vb��6tۈU��do�m]F��K�� m~Z��Y�T�v�G���I�vr����* **蠌�"*ŉFMBp��C��ާ �f�C�峪�>{TX�����:Nu��� z9�rqN?>����a�ŵX/�5B*_�U|iD� k�!�� �BrGAt�@(M���%�K�FP�,�ً�˃�.����r7v=ޅ;?����.fx��� ƶ�0�5�?,V���n�:�H��`��8v�<2J���H��BI]-j	e�梲�� Q ��0���9IŖ'�g"$*yť�.,Fe]#_�*��:JNh��N'%�&c��z׬Ã�/#3%R�"59Y��:>>At��*k���Ŋ�~���C��~�b�g��и\LL����3�I�j��0�y6��0�+XA���G a�.S|�M �$��b�G\=��n�ǡu(���W�?�MpR���x�Lxό�zf:�cCW�\���F�99��ww@������A䋤����td��s�3�)�KG�O�Ր>>�w ��V��ح��
tJ"��r{Q@�!��k� !��u�ȫ'T�J�'AT�φ�v1($h7�>�U9��'&�)�OmΧ��@�@� �
��|�?��IU܂Q�.Z�����,@3�̧<S3<4!���\o��� )��|Bh�R@�"��Ȟ���P����sB 6�9y��?���k/�E��'� t,��`E�ɜΓ9�F���,��U���xD!���S�Q`��FBV���'8`���LƠ�0Y���L6��p�\�e�1vKN��hCp�	��c&�
>Oq��)6�ʌt1B;m��s\�<��@�Hp�D���_@�Y�H�h�_M���	���Yn/C��@�f�K�&�h���=�_Y�<��1�[����1�Z�J:g��E! 5��0�|���9�)���U%�+K���Ū�T���'�<�~�S|����y�"�܋S��O�Ǖ;����0���Y�\:m���*��υ.MP��@�)�^	�T�Pc��;�*�Ϛ�N���M���4��ǔ�(S�J�W�s(��y���R��gV� :���1i������4�G�BU��A�dƹ� ���)�1�@�%�{9���
Ǝ�
4%��a�>--�ae��PU}��&R4�& *ݎL�N #x��l$T 1-%E�=)�r�L�rp>e���Mk��(�(�6
o��
		�
�j�5j���NQy��'���RTN���J�g�tf@���:i
U�l	4J�(�q�RQ;e��o��Bs4L%T�wE1 �0���1��5
��?�[���*�
�8-&�,�@������k׆�
dk�˺r���k��D=�*����j�T�)��~����+��ǀFer����xZ�S�X�*�XV����;;�ZJްƹڱ�G���:�}�t����5\��B��:���|�`̶=�cBfvЏq�q��x�8�����f�������ձ𞟋���*�S��Mq(&6&í!I��Q*��4�p�p��Ý�Wq��8t�V��Ō�%��i5n�Ah]ܳ"1�o^�����_���ݸ�������a�3��φU�+|J"������������|�?�ů>D���0
�;9����Cϛ0�qQ�X����ӯ���w|��oq�7p��{�r�$<�����kg�h�� T�>
FR����Վ�ϖ;����~�~�C���0m��|U�iYKCa@�ԏ���5�p��x��+�����wb|�;}�`��P��8�=2罷��S!�����k.@��R��AiWJ�k1c�|�]ۀ5�|�>���Z4��Ђ�u*��l�,TJg�[���0�nk]�s���O��5����5��-��[�!&��0�ׁ��&�:c5�)�`6�
�����)F���]��t�0��r��u�~�$�x�e�e�
�^v��� ������UN�е5ܦZYٺ:���C!aU��;-�<��@%
������>��VXگ�(��J�m�zT�,Rw��Ū� ��.�����|t�h�>V+ � �BC�W9�Vʧ��,[t|�Z.qE�J�O��1����%'t���݆ï���w�`����M�G�'"�_����8�V䢬��6ay;�h�|�[0Guox�����KJ�������������'��ǟb��-زc'�<�>��C�p�2��X�b9��{_~��>�X�
`���C;}[�ϑ�p��u;uZ)�'Μ���p��Y>v
#�.*������?�o��;���{ؾw;��Z�Y-Mh\6e�+�^�M��zv<�15����A�B6v���Ǟ���Gǰ��l}r��F��u*�v�`�`�Lk=�F���R S��*w4WL�-i{
�
>	��§Z�۴�
�@�����-�wbÅ�?�� �A��:1o�r4�kFU�LU�Z�E�Ѕ���s���*����:���.$��ط��`����T+�6�^B�PZ�y¦@�!������(�.(�� ��� ��݉C��b!e�p;p� ��4���FCq��ϧ
�s tE�_Yu���9���=J�[s��?��7��jU	��Z��^��`3�%3X����c3'G蘛aZHn<z��7�#0&�|���×�46����BD%$a��7�J�p����k��5Ӧ�ceG���J����- �敡��	�Ʌ�����G8&���9	�����ؿ��oz�35%�1Q��%���b_�7��
�%u(�����b��C�Ds��)�Q��,S�h`t��	�!��N�$�@���L�%��A t:O򇽋7����p$�faeg7�{��Y\W�)l�� ڛB�ؙ����x�Ug�re=�iú�;�}i���~+!���]�`s���* �@�F%P
t򷒜��4�{��Е^5ET�T�S�S)�_:������`dׇ �1yu��:�4��P�
m%[B���*��|* %djATL�S�RQ9e���Jn�@�@�,��K8O�>�ܮH�s%�(@�~@E���DZ��	��t�r��J�����6��#;��p��Gϑ=�������˸x��l�CPY2���a���YX���N�~��	=Nea�����`�� ����:�1��L�1h�2�+SU	��@6�Y��W�BǏ�gK�$��$������F������N���jK�<-�I;C;K���M��]⶗i2�D0�Dp|�. �:�o�L��"��@��'M�Şnof�˦>c��L-LpA ����t͹�a�v�&Ŋ�	��Mu��X��[�fb.&Gc����N�e���s�~��O����~�N���޷}�&��W6@F�aD ��[�� �3��7�j�U�z���!x�	|j�O��e]>��~���3�U����8����M󳇎���:A?p�f��=�������\�Ć�������k�s���v������%��U���k+�	�[)
���I��4)$�8U�UM�F$M H F�G���h`�_�ȑ|Q�2*���(��b2.������k�U-Y�*�J��D��R����CY TBoe���ee##5E��
`Jx���R�V��r\Bo@�]�Hح��$�I��̛�6��;A�#���n�ע�A�d	/���Vj[p	/���0��Zp�k��(��P�p�����rQAE��,�(�RT����G���r|���(�US�+����(�Z��U��ʴRW�&b
G��U�Ӈ�.j���ke3k�� t����n�a�`kg[8x8�a:����8ɂ`fL3��>O��`f�HG�Ǻ�2aL�'�(a
�R<a���?^��꭪ފ�)9��<P�	�:�ʣ`��w���AnN�ƥ��p��Y�z�6�>�ݗ�~�l�X��?y�����w��[���?ǝ��`�i:���c�~��ʁI�D8f��zh!�^؍�'����?�ǿ�)~��pkO��]���a�2��w/a��U\{�!>�ŏ��/���'���Kh��Eث���Ø�^C4�Ί����3f{��6�`�7��_����7x���1�g%�'C_�U �to�U=�����O������{6br4�)�v�J�R��^��0�%{����wF:b#��Hh��Z��(Gо��qyP �~,|ZW��𙿾E��Q��s-G��
M���L�����[b#���4���:l�t��M" �7���3��!Q��OC>!v��l���Ŷ������<�������b����6�0Y�Rh�@-�j���[Q?@��*T���"����R%W�SBo���J(��V-(�1�аs����(��F��$xv�$���b������CU�eg�K�/k=)J�;F�9F�$lJ�����p��>§ "�[�L��	A-2�M���u����,}���7`�㣸�����-����ipuŔ(�& �,s����]�q����t{����p��]����9r�4�O�����ؼu6mَW^}��_G��u8:2��K�T�ۖU+Q�4�V����x����r��'ϞWo%�S*�ʼ��n�W0r��I�p��_������˯��|������o�7?~;�ƂU-��|>f.����*d6�>��F?;�Sc}����t�?Q>�\0�o!��4����vc���轳��uk���<M(<�s���[�E����
0@��2��T�sT9Ղ�_ ��~|�on���F�UUpo��֫{18�U���.�ۉ�[��~h>*�; ݧP)j� ���{bў��W�{��@���!)Dtu-V񁓾@��i�R���NUt������S��:ݭ���#�����K받���B?��Wz�{CBp��F�\�,|>/��y *a����Nt�%���:�zuN~0�%����҇�§>4cX�Y�f���) ���������f,\H�KGrv���������kiErf���x�b�����?�+~��?`�ÈMNÅ��շ�P�ݖT�"15�e�(.i@@@[:@	�4a:
s+нf -�#:<���'�F"%=�q��)*"���a.�#������D$�"8V@3�~Q��th	R򪐜W���b�'d�nW�xa� �*���Oܽ#0~�?	�.��ؐ����1�(��G�iq����0�vn0�3���j,LL���e����ŅM�p{���7�o*9	���"�J56O-t*�<	��s5?�k.u+��>��k�1�Q�<:W�%�PQC��X��f��-9s#�?+y�R�(X)���M=� Y��MM�[�E�I�`���
DG!�Y�qY&ʨ��
�����@����D+8^��@s��+*a��>HՓN�w
��F�d:5i%Q� ���d����o<&�����/��*.=��%C혖��,���23 �Y0L!,$O�I^ ʤ+�8D>�m��m��qz���ل�VK�YY`%��fS�����f#}t���NW��1�6p�":l�� tx@>�px� zV��y�v�v�pz�ۉ]�Z�B`��]#�\�4�/v�`)��J.?c��¦�w��gM��:
�DM���e��[S\�5�+#U��9��r��`�xs���S��j�R�t�D��4ԇ?~�	~��W������ۯ@c}_'Ο:��7��(�d�6D)^0����*6$E�F���1��~�J���bR�H�ϥ���ۗgBo%7U�ou�RxH?�S9�:��挩|����Cq[R�"�.�阔 ��	0�&x�8����j�i�揨�$�,oE�`�R3��4U�i��maC�G�Ђ��1_{Bj�����.�4�t8i�5M�!E���$ �H��"Q4%\W�L�7��/{2���b;UX�(vr-|
D	�*�-2$UnF���I.;���[��Jhr|���\m����r=���LW�:9a�������Ըl*QS�h&ʤ�^��|N	���?��G�1]1��E���Mާ����e[�"��̗qɛ�S�h8�qQ����}�ta���s�����_�F�R�r/e[	��U�ABv�4���ʺRdJr@%�666Vu�b���T��X����V��$G��~9�r�%�c5��VJCތbd6��Cbu:r�"uV
BJ�,fzcr�&��a��S�/2���D�g�3t�]U!"�E�d�S�>E	�<PQB*�`W
[~��	�MY�rn'��v����p�����c���Kx�{���E��:���	޾��/���K���W#���SQ��5�B!�C�dB|m���Ń��_���>��7��?��	�ß�����s�G������|�!n��
6_F��B��y�*�1�Q0�ÙqJ5c[f��cL�Z��g�������7_`��N�Dy� e:�J�aVc	������%x��������Op��0�2"��a��)p�1=D9��2���4����K�Q�^��.]O�6�F�A�}X0
��~�k�R<�$�V�@� �LWm��ؙ�Лh� T
�(E�@��;��[�3�%Ѩ霁��[p�����G���=|���|[^9�����'��������%hܳ ���r+�Ox�\�"	��TJf��Y*�V�	|J8� ��n�PJ,���	�TL T��fw+SJhw	r�
���>C�C��r���+�����������"�
@i-����oR}|��Q�����C���,ikC���U�F�� �64wɩv����؋�-$Զ��D��nN��8����}+��?���_R�Znk��'�.������h����y&��Í{���ۯ���^�����O����@�@?�����q	�X�a3<zY��nܱw��z髒%6m���K�zh �GN������]ܺ� �O�Ů�p��I\�}/<z��7n��O��I(=��z�C|������w���	�%�ܸ���cQ�r�Z��}Q=��s�R��ؒD��D�f�A�t�w����1ՁM�3�-ƙ�n`���X��^lr�@��A,>�����`d�q)Ar1�oU@) �r6	�bZ�SBl�`�PQL��s�UE�@�k t��Ř}�}@�X6�n?ޡ��n��C�����к��і��[;=��y��
>.B����$�t>���{[Ѿg1��^�����Xg�P�EBp;�t}����
���� �gL{��ki�9���@�_��o�b͵n�K"P��E�>t�!z�J"�m?+!��D��n�՟^���;�6/S�\`5A涺��:��vV���c�� {:�M��a���q��((DYM�.Em�,��hBۚn$e�`��Dx��~�|�o܂�'Fp��iV�@*���3�/D�)�iDZfb�� ?�hs���٘Y: "$
��R�? aa���E�" 4S�<QXY����U�[ϠxD��#����u�
U�( :�E5����\�O �BjN	b��!Ň��#����kd�xF>��<1���}�y.i��ݺ��e����G6���
@m-1�\.~nș�I�\��������x�S ]J ]~��x���(�ʇS�ۦ�'`yV��1�|�^P*j�2��FS�pG�O�����!*\�hN]rF�a�"D9���.UpE�̭�(�bZ����Y�Tk�xJ���J��z�
Vk4�*P+ Zʆ�LT�Z�, ���OP�������Ȣc�'��r�U����H�D	�-
Qݰ�&V� }f:�
#a�B�>]w�O?�CB襇��rS7|
b`��K6䖙�����K�Ռ�
@m5�x�ф娘	H��C��!j�T�Vs#��ڌ�����MU��s��b��VXa��v9�b����+ӱ8���R�)y�z8�y�	�bF�2���'���:M�W�g���p�����5��Z�@y��H�%��%#�WL�
8Mp�{&�]�4S&
�e�\Kܲ����ָ�����9N٘���Z��{#��]��hw4�,K#��� ��o�:��g��?��ｉ�7����cxt�:~��G8q|\}ݠ?�6�0N�C�p�
�����1�19�nT��Ϟf8ZxH
#�������+�����C�Q�b~�^���s}�6��{)��R�έF��n�l��u�ϟc�p���������3��o���3g��p,a��6e"�;;���vN�q��GK+s����f��:��M�
�h<t4�(!�>
&�bb�:;F�L�Jr<2�*�F�� ��(0 ��O!�Y�3�V�J ML�%y�S&LT
��������^	#�Je\���PS���U:E��5ɴ��ts7gUlH;>�& *�-���*!��;M)��~5�Evvt"|�-��Lۧ�(���zbn�v%��=���{$0)��:�h	|j`��V;�Z���r�d\�I��1�US Y�_ʹ�>��k�Q Us	�<�(��~�g0�o��$�jbi;gPg�~�������f��'�&f�# �����U��gd6݊���hX�y�� �)	ш*�BPa8ܒ���	]o[�L��Բ8L���
I����>��)}��@%WBpǕG���m~ ܋"�x��zt��é{ø��^x�2�=:���>{���������M\}�
N�����0�G®Y��*Ca�6ˬ<\U�o|��zt�ޅ㏯���������?��o���|������_��o��?�
o}���]���H\T����,?XK�-l�:u�����5%��\�B�x�?���?��o�x�?���=�MOB�/�	����0M�y�,X׎���_��O��Ͼ�ٻY���i�0X�	��p�Q �iHE��<�B@�VU=���I�����hBpE�~@�v�Vp�r(J�����nL�q�8�L0���#<�r0�g>V����{q�-�ko��;#8��i�|�zonT!��#�@�@Áf�����P�o.f�]�{�Q�s*T�i�R.U�[BfqJ�jP�cf옧���S�o%T*��)��J\�/�Pr@�@eX����V}
����\��ڭ���m;�����U���J�+R��U��J.�(��&��! �� �s]���=J�\xl�R?<e����J��B�b�{-���z�	?-�f޷E�����#��߽�����Q� �t@e[�2C����<�.����[���^9vw_�����gx��������f/[�]=�(-�B��.4�,Ɗ�58�Vtv�f�Lt�ź�۱�����®��y�}���FET��w����ʤ��W_��o���?������?���O�����_���k�~h?�6bA�2T,jD�R$�d � �E1�C`Z0�>���6�������ߋo]Î�'�{76�r��:�BoWH��n޿v4�Y�{���Hx;N(H�|�N1��/�E���P��@e�TI[���#|&���;���>l��Cg��gx� ��^�9���P��������& ���h�:K�n�s�R�PM��� ��)�@�
n���>݁�#��l��fEv���>xv?��s���'|���F�q������ ����j�\�T��P\-�>�|�nXh�� �R�h��ҭ�Ё�|V_�!���㒦��G{p��$̄W`j�3������lm�agg;{:<�������V��^�����))CVaf̙��;w�p�jꑔ�����8͋ *����9�����u�(.[���l��a._���(��%�r?���i	|	�!!�HJ�AlT
}6ܞ��D�ƋQ0��� BC	�����**ƶ}�Q?w1�M���W"�s�U��PP�����|w ��n�!��F�,żVB��~�_�y%�N�#��n#1�#�^1<V:����F8�CfQ	f/nE}�\x�`�DG{,��`Ic�ˉ�Ho�C��zԭ���K��}y-V���hQ�Wc�	�%8�B� ��~j�P͸�%{�e�?!T�~���D5E�V��)�S�T�s��64ʎ,�CNc��BQ� ��	63��g*�xZ�V��'�Rf��sV"��1Y�H�vEJ�$�։*�ꨄ��BJؓ�B���/�CAY�F!4������|?�Oh:��V��)D��#��R��y9�����x������ǋﾆ3w�`��Lˍ�a�d��i��Bpͳ�U_�ބ�'MD�%1��A�ȝl�J+}̵6�B��XE��25G��9��`�	�2.��a��%vX��sC5��q.;I��"C� z�@za�.r���1H}\7�Ǎ�F���� p�|��]~M ��)v��z�h,.s����7�ʴ�:�����W��q���\q��7\�p��
#��p������� �'�b;t��	jֱ���n���e�7?�Ͼ��|�)�p����7?��<�����Ê��}�/Lҽ���߂p�< �DzE4>#
K�3U���B�j�=k�>����P�OKLP=�jz��ѧ]�>U��P�4U�VW��x�4q2k�c	4���U3+Ѽd�+дp��;�������O������x��W������?���x�6l� �Y�,�Ȗd13[��L�eff33�c�3c3%3��f�L��nv�I6���_��ꉓ�|�����}�GUWWUWWWw=��p��i��f&$�����N�N�s$��m��L��yc#X��O�������"x���@G[�S2iR�V��	q�c!i*UU%�'\M�o��N�3�����d[	��U�%8����=�JRA��~+�}F�G �x�y���R�V��J�M����zBڂ��
�Ĩdt%ӹ`�<U=7&"��Q�i���	:��EU�MaM�,�)x�c���5�]5�4"	FYW޷꜈�)�9՞�����6Ҧ3��G����Z����#�_ٟf�{ϝT��TUgooBTڞNAT >5�s+�-�Ș�r^��d���K�['�����{vrv�����1� u�p����IH�:b��"b�0<:��%�X�u^y�1~�o?����[n���C&Z0�����|d�� 23~�>�G|Z:�"����x��j�r�H;gi�7�!0��ol^�K#�Ԕa���P8V��.�� ?�X���}�|��O�Χ/�������������ǟ��eO��W�����5�7#�!��?X@�h��C��{�qC�kb�:A0�j�5���f���O����o����Gￊ�/����y��>œ/�Ʈ�'Z����W��{�iH�U�)�ӛc�S�ڀ������iQ�Ɩ�_��q��M�z�!*&a������H�|��y�,���ר�럽�g���/�AFc1f��aF�#�Nۢ0U�2��~
�����#i�'�����؂�,k.cyQ *=�6�S���2�D�vtK=����z�"��+���:l�} �����������QB`?־�������憃݌N��{�P��	uZQ���ь���h;�u��-(�ք�xS-�6�*X��c�ȝ(C��F4�hS!=�
4K�Pm&TD5UrT���
��SUqK��P�/O᳔ -��ț,"r[4��./��9tI��	>��ӃDG?:��v���L��u�9�TU���pG�L�O�j����j���	ρ3��Y)���7����<5���7V���YD�p�,���YE����-#F�u�>��W~�6|�):7�%�ihZ�m#=�ܶ[wn���1L��@K[+������m혜\����b|b-F�.�ֽ��~�VV�#�� }K�`1�ٿr��|>z�M\~�"��s��5��2����ѷ?�k＋w?�?��_����g�	P�o�#>���x���8�:4�]>���NT���Y���lDT$!�4A9��K�w�}�k5]e>�X.�|q�x;_>�U�wa�뇱��^��ݢ�N!����D��Qt^\�����P/ڏtĢ R[�V��`��p���z�Oϋ��%���v��ʀjJ�����7��C=���\��w	��{���N�>��/�nP����7��v��>t�{��kK�sy��.����C�xaD �k_�@ln�z��� ]�`��ߊ5�/n�����V��ft:��3��U�C!�Ւ���o����`xa�t���	�?��c5c���Jl=�Je@w���ƚ��|�u��Vc��c�/cD:��ǜ\ች�z���T54z��D����+�0 �6��
1z�S8���h�Dp�7�x�@�R�f�`����)�8�����`�_V��c�DCJ�jP^W����uw�yQ;2�s�0;��������?(��E^1�&�����ؼur�QVQ���n�,�EZv!�o٭.����������/0�7n��;���y�yK'����Eddbbc�T|,F�1�/E��M�C^E#ZπHx�G .� ujq];|B��4?��,�,AZN	q�ck������L�>�1oA4��c���ȸ<DDg��#��f4	�h!�3K����+�m�?[Ӎ�A�Ө�X��U�|y��������$3-���R~,�'ܡ�ģĹ%�������D��]ye�M�*|��N�1����E��Q�"Ym�ȩ�@�EU�(��M>�!s%�L�)�#Q� "s��,o�9����Ȫ�����}L�儘l��,
��	(lJD~c,�]�a���-C��S���/�A�U#�����.��4��Coę,Ȥr� i��H����H$�'���7�PxdG�ir{/�ƍ'�q��ѵ��i��L] �� 3e��� �Gc~c:��p�~�YpJ)�bA���Q���g��($>W�a��L��؈�s:h�����)��8��26�)�Y��?u�ᢞ�p;S�"ÝH\�e\%4��������q���p�qO��B�3��.���!�j�x��}�xɄ˸������.1|[eV�������q�q�\���p�� ��Lp����m�^�v�]'\�6�is=��#V���Z��M�g�=�x��^��g� � �rw�O���~�9�}�>��-����ݺ�KWN����mf�8��	�a���\6#���'�$�H���@�D�a���Nl�(%�b�tĩN5�YŘ���p>fTH�����,�s�2Ne^�����|���PL�ry��e3��\�7�e���t2�cZ�`t>tR]1-݃�y�NĂ/xx���y6�0�ߗ�T4חct�۷m¹sg��g�u^�u�᏿Ï��X2:��R]���A�~�	�nn������v603��U/�R����Y��T��H�N@*��� S�xj;�l
�X2��F�8MUT-"�� �Z��\H0)�	IFS�R�V�{m �TX�"�4�5�2�C9�dl)|-9V�EV2��� A� �޼�D�!)!Iq����R�꺂Mɘ�T�6�Cͻg���_��ג㑩��+�d-V�nn��??oB݅��Յ�t�l+�L2���&]��bg'[��H��=�L�\>�l��WɆ
"�3�s-���|8�����F��t���dg�ގ���Ē����2h ϭ�=׵��j�F0�0���.��?!�<�A���4��ɕx�՗p��E|����Ϳ�
������}�w����Eo5�J��0W�KGp�܂x�-�GBq2\=�7~���:��i�����h�=t"]a�G�:�Q0Ϗ�`����0�9�0X8���������wq��I��{go��s{����80�}�^��wn�d�	.0��͹%V��h  =@¿r�b�P��Ebv]4L
�a��؁�X�ѓкu���Ѷn1�L�m�(j����Q������O0�¹i!��aٕ���j��_OOz�m�T38?���i����$��p���e����XUDA7�C�!�g�$^��#<��M���۸*��/¬ G�z�$�ف�Ṛͩd@����Dv�"i��K+Q<^����l�ª�U���laW��	����
+oH�7,,U�G�YN`����~�k��˱�D�T�m<؃�}�Ğ6��,�ވ���=jw7�nO������ۂ:��� ��ن�M��Z�lJ�|�P:R��5[�и���jQ����L7�vs#�67�vS�z\M�Vo�G�V��˺E�e(�(G�dS'+�c	�/[W��MU�%@�y��`��1,&d�,gy��9;��S�h9��)�����<oDi��Bd},�����2���?v}=V�ތQ���O-#<����<��?L\��\�����FYƓ�z���3,����#�:Y�ﹰR}c��c��zl|�G?���?~������Q��=놱��Fl8�vm��M����W���˼�����	9iy�X>�o��m����X�bDuT\Y���<��W�������'p��=\�}W���+O_�����{}����W����������;�;�Y���}<y�1'�br���n�U]��o)Fjm&k�S�����3a�aX�{o'�X̀��
*������:�=;���a�;G���F,�1��CW��,ϑ�T|~D���s�����~�����$�e,P�HI�=%8]6K���g�E'��-�91�6�S��)M�N��8��cD��^�Ŧk�0yfƎ�Ǫ�U��ݣh�ҧ��j ���M;:в{Z�v�m�&�1�g]Ɇ�E������V��{g�7T�е�Z
}=1���1Bq�4apr)��k.q{A�� �6�c�*NWaB�y��$@'xNr* ]���(/\-@W+��Qu��j�+UC�ŌA"��2?~H���z���<@�.KUϕ�BL7K1~w.��:N~t�8�ǂ4WX���� 5���l;Xؘ���机�w#4{�=8���x,��FAY)���}mX�ؔx��Cx\$"���ÂyX������������v�'BϠ��5�����3����w���X�~"��0o�TW
F����D�us��2����G#*:�,��_���J��g1�r9�҈�|��w 9�A1���H B�/켠(���Wp�j��� �Fz^9���� مu(*oED�D!:!3���je�	��H�n�_t���`�b�Y6z��Lu��K���v�#�WbË;���Z@��)��]�(<�8U ��}
�
�����C�\WV�T�Ӿ�M}�Ymqȕ��T汐p鍶P�+#��(Z�Juܼ*�PZ#𔪻|�5�2��0X�̪��7���L��3�/s8�Zb^�Bz"N��aaQ0
�Pٚ���dM�]�H�WC�V� �<�|�x�7�Uq\C�Fa!ySN%C�D�&5$7y�p'��/@ْn�xw^}�[O?�f!.�Z��BP0�e�@������PU��������(_Մ�����@^��l�QF�5��c�,,64ƨ��`�@�&@�mz:�6���^47�q��������Y:*z���&�)|^1��k���v�/
��_��u�p���3�əD�&�/��x$Sn����L�����a�5������^"<�,�`�	�ۘ⁽�����7;���[,�^��-�q���a�'z�7�S�~X�j�v�~��,d�������9��Wpx�ٻ�N�@�;j[+��=wS���U�n�k�����S����>�R�U ZD|Jp~���IxjC*��t�Ǽ�g�ڝQ9�PBS2��Q-�,'Q*�kS��������56�����F��f��0�0���n�5 ��l�4�:���I�6�&����ߥh�����ȋ
DUf"����^ڳ����}�y�^|({?�KO◿�9��7��ʱQX�vs�Λ��|ɮ9D�pw�ԙ �� jfb���
b|�|���I�i���2A�d?%'xp
t<�ɸIN�-�M� JO��*���|>���؈(B0� �S�|zIgC��:9��v$��^+M�Z+�U�O��c����a�"
��
ވn�(H��J��Ym/h���ڭ��+��,��4��kt%��yMɤ�{�e��,)��*mK��Pw>��??���?�B7��h�l/�V�� ��w#@�%)YVyO|n� �U�P�j��JU���Y�c��s��S���-��禲�<���Z��9���/ω���[ �����,--`ff� ��h/ow� **�!����ā};������'������y���O���c�c���X�z UM��,JD\Z��}��cߘZ3���n�Ʈ�б1�m�7�+s��MF�ì8/�.��su*lJ㉺��9E��/���m�"�P��l1�-�g$֦ �<V�4?�g�c^Q|k`W��������HX�G��.3�B1�S���5F���Y�Gú*��0�����<�xH4]��p�<L�wǴ$O�,�"øM"lZS1�#V�a;��@�Mö$5�>V��6Ĩ��Tm��`&�3���0��~iLʉt���874m_��>}/}�����DR]!�"=a���![zÜ��"��
n*Ϩ�<$� }��+�PL���+ΌcA4p� �:�Q��X@o?܏.Bt���ѐd�%�X&`a��X��O0�B�A�u:Q��U��P�莆�5S�'<�����Z�߸�]��*��^l�UGC�E�`r^�����$2+��(��q�a����*!�eh�x9J'*P����o�Aʐe����RT�jD���X"�o� �5�L��A�
<�6],7��E���@�((�y��6�}�GUK[���-�� �re�>��y��K��
�K$�'e�_��!bY��h#���?��ے+����
��^>��_������o��/���;'q��9�~��=~	�����	�|�:�;����V�c��ص{�oZ��7`t��m�K8m�jAEsz�`Ӂm8s����{�ſ�3~��?ⷿ�~�/�ƿ��w�����;��������vp+V�����#�h��g�V��f�!�U�+KBly"���k�'�e,_7���vƳ��Ѻ�����.a�ۧ���������Xrs\%�$�RM����cyX����'�x>5Uo��O	��7����&d�P��f��g���z*���� ��:G�-�֛;���F�:�����N�zv/U �h�:�nhE��v4�$>��ܶm':v��P��"�S��v����1��K��c��躇�U(�������� ]yy�'X�g,S��K ��@oL�^LWb	������Ā|�.��uq�_�S����׽�� ���O�!�+�	�0v�#�i0cAS jeg[�90��@@X ^8q��'������DT������w~�=T�U�7��㉷h�`��\��&����+q��Ҋz~9vb톭���Ks+ڻ04�
�e5#<�2PRZ���8ތ��S2�p��9�-���\�-�Į�{���Q��i�+��ۼ�^FTr�������Z�UM�)�Cqm+
���Y\�Լ2��R72!���J�W@�r%)��+�w����E$@�g\['o���ar�6�ٹ��`����#AoBF�|҃\QO)�'[y���p�:ǒ˫�p�/��3�r=���p��F��D�<d��*��_W}��@�y��%Fsy��[��I���g��O|�7ơ�1�E�e8,\g��{��LTX���v�	!n��v��sF8��Q(nJe$�ȯ#0�Z�!Ȫ�|҈��3�&Q�BhY4 �y�Hb�%� Xe@����N,�ŹÂ���Ÿ������������u��e3BǘX0$0L	����� Շ7�U���u4��B`�<,��B6?���F(!ؚ̍�ij�.�Y�ҝ��^�6��"��_���\B�m�c��6f8Bܝ 8O�����g����
�ay���I�
��Ƈ�AR���L����x���>g�x$a8�%��5a��GɊ�dJd2�s���5��C�K#���/Y�%[S�do�GN6x��Gx��{D�U�\�!@�q�Z�f�c'�\���.@?���s�@����E���.����v� Nه/^���)o`+�L �,��`��Ba������@�8�S ���8���Pf�Ih� &g>�q�ȘU���WEa&�c�T�`�t�d:��1-ǟ�$6���Ȓ���3�0#����_�?f�{C/atc�q���Pر@=�8��a�cX�`���X?�E�!S�����d�����+p��!\�|	=��W�֋����>ǿ��7L���N�ֈ
�?�7���\{�Ӊ(q���5,�
����F )��I�-�Gb\�nD��J�XM�C@��Om�[A�&�i�(p���B*A�����zj�s�q{Vŋ0Z��x?��+��j�)�H�H��@U��l��d�OɊ
>�9���W *�%�s��w����s]�;`�)�e����C�H�\A���\�ͅ�#�Y��kh��N�d�E��>/pTmL]��΀���|�ؤd��7��/��T �ELz�n|���!2��U�g ���y`.-�����ڐ���Mm�Y����$��y�V�j�2ƨ,�v�A|�� �v�,,M�P#8:�"(�Qѡ���T 5�5�]m����e���������:~?o�(ä��=~&6-AM[�%@b|���� ���a^��[�b����sъ!�|��� ��N���H	�Uv8�3��K�YD©4Ε��Kh��%ý6	NE�L��(gX&��*���sa��Ht�Y�|�J�����0��w�2sZ�`T��P�3f4z-���:����2��(����>{aF�L��aZ�¸*F����@���-�0nOVY�Y�	0Z���̯�)ؔ��X$4���T��WGà$��2�?|�~6����%�
���>�%v+�������p���8y�2�
`=�~�=��o�|ޟ|`���� �Ȯ|�� y�K�P�����Շ�ǰ���C�V� ��G��BZT�����<ԏ΃}h�T��'6+w���ؔ�v��ϊ�-�g��ۉο��D(����d�|����ڬ:��Z���*R�V��\C$�q�d87h2�2/�h*�r^�P��L�Dg� t����
e���ue��ݤzO]vsB�TPb����G����k+�}~1���0܆�e�ǇXn_���ȥ	�l.mm��ي]O_��;Y�Sп�t���
��,�K&���d�!��;���3D���\��Y�[v}�/n��[���6�zG^=��O��·��҇O��������Ϝy������ƅ3�q��i���)nݻ�=/������l�*,[ǲ�ITw4�,W�Ɓ6,^��oǹ�q�͗���o�ݏ��ӷ��ƃ�8u�$�߁��+�:Ԍ��"���E��G�j��bUK����Pf�Kڊ�:�Bڊ�`��bJ1vt-��z�����Naǳ�����E��#M����4�9,0�Āx最S���h�N���)�O�3� =IxJL�SB�{bH�s��x{F���=9��^܇u�`�Q��V,%D{�,S �^ӆ���Z'�p�w�{�U�VT��m�!TuHt�]{�п�#������o���v�P���ħd@��٤ :B]K��������2���EG!T��d@�//C���/���S��0��K�Ѕ嘸�'?=��g#�!\u@d`��ٺ0�6 @-a�0s�:������l�~p���Aa9і��Қ
;{_}�B����ؔ�D��o>�#B�������B�8|	Ɇ�.�=p=�QUۈ�żЖ�DCkJ*�1<:���!+�>��,D�ۋ��1�����M��E�8s�<z��������`�����{v�˱ 4M]��n����:��q�w ���ټ�U"��JuB��]�𸅘�G7_X�{��=�+U[���T"7	!ᙘ���D��&�'$
��G��_���Z�����y���5L��&:0�k�����-�=7iS���B��UD�' ��2t�%�J�?�ܾ��b��iAɲ�)�F��� %0@�Nha%�)�	�<>��+�F!�7鼺"T���x�v�X+WC�9���֮s�3�1�����`���N�g!#l�
��ɂ@n]<
��P�N��&q���XdU�#�:Y�	�i<2Kc�^Dt�#� 	QHnN�!j��Q,^�o���~�c|��Ǩ�k��[����,��8' y��S{�׹��_]
2��а�ũ!��A�UBD6[c��|l$����F��@��4����:]�TcD�nGK�1���j���s�>g�����p�x:�2>�z-AyO�9�E��@R��>0��G��xb���eb�	s;��	�W/��e��|<�0�$�)pU�O>&d_��@���ᑃ;��	���|�D�ޙk�����9�8%l���/,p�jK4��A��N*�bK3.��X[-�N.��k�e��v5��ｏ�~�=ķ�@����ݡ�AlJ{J��*�|��Δ�
4Y�EA�-��T�M���p�I��e�0*��Iy4�+c�UZ%�X�^�B��lr?9A�������qZ�@�����F���ёA�e��8�C�����l-fA�7�������v�M�p�DTb0�R�Q���Zl(���X_��^֮^�C�����#x����g�~�>��,��/��l+X�[�=�~&s]�Ĝ���,�Mad��j+k�_�ҋ���Xr�1Pj�)���ꮂT�d�b��"I�;�\p*�e}�6"8TS���X�҉�t*$��%d^<��$��I
�!�O�[	V�p%�*� 	�T���F:_��� :%���!����m�	1ɠj{ɕ����r\._G^[0@P?_�W�u�R�;��h:2">�lf+0FD�!8DP�I�j0�2�S���"������TVT ��u���2�l��쨪�JSp)�M@��xj����J�����z�i'����T�)��KJJB(߳�������-�-L`bj G'[�?411a��
��L$'D�������ǟ��g�=����+�;s;�o��x7J곑V��L^����X?�x�C��~,[�������>r �c�h�ANg�C��싹�I�-��ua4\ʒ�\���թp�K�kM
|�x/�M�Ky,�������MUlj�`����k�	G3�Uc����~G��W�Y��̆b0�0��Nmfr��F(6G���@:�3`ڝ��T�=�0�I�a�B��A�33��1�w!t{R�ߝ��)N�x
>e*�e��k1*Uq�95"D�y�U�i<��5�Q%�$���-�sE�h3��&����}�e��}	���0u�q���`�����"��.�7�OhtO>����
��A��t���	�	N	�V;�h=ҏ��^x5m���X�x�Y(n`��~�"T�5S���٪Bz��|n�h@�߉J�T�)!�[>%j��t&Ddr*(�q=����U�d�Ui��:4p�ƭ-��h��Z�rɄJTe?WW)�~@�֗�� ��ӌ���^\~E �u9���dt��lљ!�Y�����I,�LH�l���Z,�����W�\Knz��76`�e��3,{���<�:Ih�Ю3KUT *���m	��D��㲘Ƿ���U��c��F��Co\ۂ�w��ʻ���Ç��OH������o��_�����?��j��.����+��+6�������!�4�e��u��h[�m+x�Ԡ����,�v����-�Dg1*:�Q�[��.^s-����BNcR+�W����NS��p��C�a�f]g]�y�#�8�ۇq�S8����ҁ7�c�뇱^�yw=V�(���� ˮÒh�6N���g��g����R�Ik�y>�P��߫��qB�)!�#*����:2��|6��]rl�^:�MWv`���;�I�ڳG�mC��ZT��?���� ��߃���h��2� ��f��e����^��#{{1y�� tã�_#t���XO�J�ɛT�e���[��������D�[D�^��T+��~�I��_�E�P->����l��!rk��N~r���!����9е�!�a�¦�=�h{�������Ӂ#�O�d1�3�T��e!� -]-�,�"�����($�'b�j�hl)9�!�����XHXnغ�lGS;;z�x�8������}#��E^^b��Et�x� ��|(��ӑ��P�/  DEN^!2sr��@�.FaU�ܼ�����2l��^~�C�X���Ib����h�A��r�����f�]`�H8{#(b!���\H�.��g$\=#��W��Vħ碸��7�AS_;�R#U/�Ps3�t��tD�Ģn��[yA���<W��Y5�|�� *��^^�%��|�%J���jF�R@��PLL�����h��T���e�LЂ�H�k��>�|Ʉ�š�)	�,������f_���1�F�p6��\#���D����X�-��I,�g�#�$�5q( (K;2���4Y�hM"rj��#%SJ"S���($	@	QK"A/�Y��8|�����AEg,�\a��#��͊B`���#�% ��g!&v.�:�-�AS�,�E-�VE�x8b��m�ƨ3��:��h��A��B|�q����"q��l���z8I<�#"/��&:�b:���F|N�M.�E��a�7��i��x�ţ$C Jt���g�3����x�xJ�>�����sC��@����#<��zl! %N�2�/�/���e'�{smq��<cc���f8At�1��9&��`�In7�c�$�;x܋�MQkb��ٖ�NŶQ��������1!�.���������Nƌ'����d3���v�5%@���Sz�UUg��Ft�t 4�7ܩ�����$˰(��I�t�7tB`��R
�B�_J��C7O�۲�XF���R�6%10�ƌp7���cNt �K�[^�pB2���5Hh.Alc!����S�y,x{E� 61�IȎDz�
��ƒ�/j���R�߷�З������x��=��w����7`mi�W�y��5B,9ρ���makc�:264����*s���������*�Դ�΃.w��y��@T�"�t�~����9�<GzΕq/#B��2��D���ϛ�p�Si��`靕0���ڪ�PmH6T�(YPmP^O3&�7�� :���w������ڭ����S�%���Be�O٧�3"o�OɊ��kח�=�9��v��UGFMA��o���\:��Q8�m�ڭ�S��JU���` ϙC�B=��������|��8y��mMF�g@���|M�V-ɶ2l�tr$0��e?��T��G�@]�z�����6��"B}�T$�F�z2@VF2�����O��O?� ��&�y�<|���|k�L�oy;�곐^����(�&�
�� �����э8u�8�]=�[�o���۸v�N]8�Kw�c���H�)�]���R0�,��ʂk�B̭J�GC�[�0�9�3�ِg"Ծ1���mO�MK,����0��F�2�5�Q��k��n��i��j�oA���a��f������#J�:$��e#S�iЙBx�b֢$P��tpjԗ��TLo�Ǭ�D�j��~��F��Kh�9]^���=��z���:<��`��:���P�k�kJpG��<��|��?ģ��o�U� ��sa�B�f�7�������tj6��@��ݝ���"d,)WUp�	��=��?8��C��:���!4�p���m#��Dg�^��j�Ѹw�Bg��M�xVl�*�x�mkD�V	�ok���-uj��ɨ���[�U�BuSC���hU! ��ު�IFT����i�v���|
0��6T!T2�S�qk�2�
���j�� Z���e��iA?�PP�)�=���J�����S�����1���>����&�����{۱��N,���4m@�;@'��NB��0�tT2mKTЎӣh�ꢜ�v��6ta1���Ze��%0�pw�Jrmi��v�?����_��w����S���O~�c��~�?���o��w�����r�6�޹�`�04�-=Ȫ(DFy�UEȗlf[1ʻ+P=P���j������ ��������E��\Oٍ9H,KBD^љ���D��*�p����f�uу�Ls�������7N��O_��/na������j+=����i��ߞT59_À���� ����,H�Jtʼ�B�A������Ю3��7�3�A座e���=�z1z|)<:�m7�`���5���
��[6ހ��z^��h��E`���@����)�O�g��N���@�>��{��tcxO&����W�]ǋBbB��tՕժ�儣 t�E��>��+c��J�s�xѭ:;�U<�g��K1ɋq͙eX�Z�Il�E���$��CZ�/�J�s1*�p���a����Ri3�߄�a~�R�s�T�\��|o�><���u/��c�f��,�8��ְ���s�䋾e#���X��G�%!4:)Y��*��t!椩���hZ�BԶ�c��m_�e5
��1�E�GlR&:�cö]X�]�#^:�ޡ��ihGyU#�Kk@���@%���$�V#;�aq�i ��C��B�e >9A�a�njB��(�ݼ����AԴt����9E�JJg�����*�y5w!��
�a	p�a�bAP<B��[Ԉ���;�a�����,T�u����jmC}W;J���� ��������9��T�Ӿ�h^�� ���32��������
�F�C���*��w2V��*C�aT>[ɀ2T�S�Mm#Pi�ߙ���hU�x
���S: *��B	�YX��v��#��ud�bE���(nJⲅ�\ +��!0	KGKX���p�������a5�&����!L]�Qb��V�&
�s��X��k����3
Z3U�5,Dvu�ʈ���"�8фg|S
܈J�X7����zy?�<�����̍�(i��U�;,R�0cf�E®"��S�b�
Ba��Ķl\�sO����\�����e�:(`Z�����j����A��.Zf���H�	�U�mo�#s̉7\ J/��)j��kS �e:w��{f���� �J0
_hZ0��3��5s}������7N�7���	N�7L��������^c<#8_��g����ʄ�6�+v�x������U�~���}��g�q����-q����9f��qh�o��.�Mfa�jn�"�'F�:#�~(-�˧p��I�'�q��S}`�2��>��J����S��J�iz��^௪ݪ΁�'Z'�X�)=؆�,|��c�Q]^�3�X��g���9�q0N��l�9A'О�@ f��Ü��aatsY8��^Q$f�D��,f	�*�ga0 za��/I����x��{��/����+���G8z�zW/���"d�a~b(ܢ�07�#�0#I�~H񛇬 ���(�t6al��ؾ'�ť+q��Y�:u�o]�;o?��ի`mn~�~^Ď�1����"����Z+�J���R�I�pq�,�F�I�ҡ�`E3􇯪V���r�tN$Uk���_2����Ǿ�aUd?��y�
�2���T�Հ������*�ܗ`P�)8$JR��Ne$UV���h��M<��@��tS �񖌟�������~�\ٷ�S�'�O����+C�xy{��Njg{;5��L�������N*\]�s	zM�T�)Um%���s�ב������z�ߗ�T&��rN�3h
0��fy�R�XBډ
�e��V *@�������Ԏe*@u��S���2���1�x�89ρ��|� 8�We>����LK����HU�������~��x�÷p��-8�#+ѻ�-�,MFBVB��1��>���g��Z�%���~�Z�޻.��k�=ŏ~�C��?�����q��#Tt7�&x>,C�!���$B�k3@}�
�C�z�g��1n��plɂ]Gl;�`ݘK�ٶ>f�0����S���Y����Q��:* �I���!8���H�JU��x��2�`ؖ ��$��*�aؑ���qj؞�uU[i���zj3�Q-F� �>���b_{�d@k5�Y�ߗ��{cf�+
����O��'?��|�&.��"2�*0��QF� '�y���V�
@=���(�rכ���
@+�6�qK�w� ��d;�_�SC�4��B�YKX��b�dw;�$vM��y�N#�u\�B����2��:5�eU�R./#.���M�(�X���,Cʴ��)l�O��V����;�TU��p��k��TځJֳi{�_��e�,��R�V�yQ1ZBx�H�D���l҄�M�6���U ���RW�5
��s�Y^���at�}D���qK��e�V��d:F����kno�R���p����4��,�k����U
�ώcÜ�v�1�N���<!��4��g	��,��W�b��	�~�	{�>��߻��?��˟^�ٷ����3����՟�_��g��?�~�}��w����Ǹq�E���Lیʖ&�X���^,,�ABn
�f �2���Ȩ�HS�V��d3�:=H���`��"<?1e	�}g�,K�O�/���Bo�!tf�`�\=̉tBbs�	�^9��߽�߿�?���ߺ�����{�����۠��қ�L[��K0�2��E�_�^:E���T��f0J���S�~��)�j�}���:N,F��!4�0�֣�,���v�]�?���� a;���j�F/w�W�Վ�X��/��;1zp�1�!N� �N�jֶ�jm���۾�GUw�$^��[����>�?u��߹v�tўN��Œ}�?��ӯ;!����o!@�c��5X~qKN/�(/�U�tR�s蹕�
t9����
����c��Xwr)��]�'���6\��@����������_��o�A�ˤ�Itj�9$YO~��#��K����n{�$��K���@KX���jlY �u�W�z̅_L8:G�x�YEp�#2>�G�壤�	���(��bS�T'D���DM�j됙_���bDƥ�?$A��)������ܰ=���j��=���f��ա��&\C�cx��b2h"��y#�Gtd"#����(�� <:��!H��%�j1�/=���ʛwə�((�|[��N����JL�oXq��Y�c�DLR�g�#�����d4�%j<P���&"��5�(i��Գ��1�����N!���Dt^�7ZЦ-�:�kAƐ�!SO�lJ�S�PA� �/ }.�L���A^����3��p-�2���ж��+Pؓ�h���j{�|��D��ymN!4�(-��S ��=%Zڒ���4D������
��v�+^?*���D�L�La��/��,\M0{�9��Ƽ��J�ALA��Q�S���2�w�؛3���K��ai$��5P��0�
uP�8�ހ׾��Pu�����n�o�ڀJtNe\jU/�����0F(��מ��W����cغ�
���
pA���Bh�����c����3Q8]�z�P:M����h8mz�ѯ?눱��8�sp�� g��U�i�i&�����M��5��}�Yx� *Ul�� }Jh>�����\��7M����x�@�ƻ,tj�=B�]	+�km������$>��}�˞�Y�u��x���O����wx��	�+vf8�k���)��{�Ͱ��g�hz��;�#&��h籴�l��f���nȊ�G-!��A�	�Ç_���@Lw5�I���hC
e3��_��z;�Д�A|N/$:�
n9��'cFi���Hﴌ�ER�-c����揔�m������?ĖGP<���`.t��=p�q������E̦@?/�E�0+��u��
��H�����+��?��!U���_����_|��x��C�m^����e'�?1�Q�⍤�xTT� 36@^�j��\���>�\�۶m©�����=�>u'Oý��p��~T�����6���p$~�76ħ5�����ڀZZ��T�b1w8;%D��EI?�A���Ӭv�O��O2j�L�YU��ia��������+mI���E�S:|J�D2�F���yfE��R�V�)�b��Cy,YIA�d%�LD.�6e��������O��rnD����+�I�Z�gLdb�/���+�zn��S�� ���18���s�T2��)��<��S����2Ʃ���~�2�s�� t��3gD !L��s�6�|lmhe�V�y�=���R`/�Q��J&Sާ��@�5�P����*�Q���S>_���|&2��� ���VB��w��������Ŏ %ڃ|��/)>
�-M�O?y�����7��+��~�w>xWn^ľvct�zGY�j&@����3��x 4��9��7䡩��KYhZ7�=�v�ҥx�7��~�?������<y�)j:����*Bۋ���5�Ӝ�Оr��V��%s�21�-N��aۚ��DX�&��!Ý��'��)&��x"� ��&�|�M��(*(�UE����0�K�@�1K�ٚ�����FD�q��e|�.oN�C��d<��o�it�u�rfԄc:�_	��PH/��#��3܀����>� �|�6n��9]5�`�t?���
���`��ޯ�aو��SUpVV��~�X�%@;���EڛM����g=�WK|J�<�Xp�(YQ� U!S�B!*�7Ԩi��&��hQ l*�2��S���m��4}�O�zʼ�Tn�ݡ2�ĢT����d?��0)��+�2� ���
�Z�r*в�U*󩲟���n���T��y��䃍%t�X^�N�����N����H��A�.2��bBr��p��RtT�LS�1��%4Y��=9�"T�y��YN�hB �A�,:��Pm��$QJx
>��AL���w��'��+,��X��o��g{q�ݣ8�����~`l����;�SO���7p��������{�g�����p��=�=rݣ�
��+#:3�!H(HB�t.V���hD������H$T�lݚ��-C޾�%����{���w6����7S��N�'=�G� �1/����ƙ��ҷ��·o�Է�b�{G��̓��l�>َ���{���,����I�\[I��P�2]��'q.LA�N�n��ǂ�籩M�S��_2���� ��������m4Un%��ږ�U�2�����C��>�]vj�<8���a�<�#k	�qt�Z��͚N���P��A����@?����C��^�	�d>��u(���]���]��׍��^p'�����䭍*�����%��*^�� ��~a��ʄ��;��*�/WUp��� T��<>@	�~�K8]���|e/^x�0
���5v�a�: ҇��5�\`��_/$�eb:�bE�[l�B$�e`av62��8O��!�HLOALr<oVQ�H�C|Z:2ʈ�®���[ <����;�Q��#��Z���ehj�Fet�ۑ�W�!���e<�X�F� ����JB\\*�B"���D�
����
�d��xґ]T���L�V��{��݅ʆ6�t�s�J�/�e���#(2�c� (>|-w��ᐇO��	�5}<G~pp���"������8T�բ���,�:��`�\k�:�K�:��0ي�m��N,S ]vm\�S���@�p�|u����7T��OU��l�6Z\����"4� -����X��l˚����( 5���9f��b��-!j�j�h�2��Ĩ&8O��;�3�`�j���V�zZ�����X��^A(���ӜN����Em9H�KBrs*2��YJ���1�X{�|��?Ǘ_�^{	eU
��i~���iA0���h8T����� f�!��<��;Wb�@=�� >@��`Y���,	�i�%[	�:B4WW93uPj��bB���7�C��.�g����,l B�[᤭)Θ��e��e���&:�e2w�{\�P j���zJ�W͉P���,����8��T�Cܽ7�O�&���ˏ$X�����p���1�%:߶0�[���'�W�1U }��	o�s�Sb�%�9�mo��v����?���F�mk���mXn4��m0�����E<�v�~�Rx�]���^�/?������G��k�1?��ޖ0�v�^��iS����;�iS ���xzQ���D�|�1/�E0)��ii�B<�}��]��>����7�wޖ��p�5�+�c<:s�a>�%I���pw��T/��*�B��1�e����~�o����s|��������p���#��L�IFtz��B0/�)��h�+AN\��|QJ��%��8-�X�l۷o���G��՗q��;�p�,^�sϝBCu9������?���N���� jin���J�4��6T;��}�ռTmU�O�S�m*kJ`*d
�8�<�O��L�
�T���+U^�'.hJ�Sz���Z.C��cA��ʫ��[w��S��JA�`T:���c�^^���u��
���@]�@e@}�d?R����ሉ�j��J�S�+U}屼����ו,���S�(�P9��X���eH�e����jY>�����.v�
���~È� ��y��u������i�a���ȹ��ZB[W:�d�5�le*��9x�TK���N�-�hmfڏ�K�~J'D�����l��~@c"B`l0����＆?�*�ӟ�o�����Ǯ�;�x� ���������;5!1�����<�1H�OEY}��v��%X�q�܇�W.��W�?�1��_���k���g�u=��a�]؅���j�̅+��W����h�Ƽ�"�w�L��N�i�oH�m]2,k	ҦTX���IЯ��̚�S�}�3�T�W��p��
D�x��W! ��F�=PCT�^�?�._K^O� �T�a���O��� k�/�|?��=<!�/=���EU�� �Lc���es���a��Ϫ@۳ӝ��a)�E�d=7��g� ��Pۉ6h[	��]��.��*tj;R��ഁ �i��f��2֦��Y��ZM+�����N}�m%aG��sy)�/��_C�Qv��l��|
<��䘤=��[�DJ�Zh1�(�R�~+��J\��Tӝʔ
@��M �N��
�#Up�=ފe�&��KP;Oh�%8��D� Q9z�em���ç�c	���.M��|��� �[B�jS��ot#��ΓK���@{���3�(�G��C�ư��j,������XzY�[M`�yVߚ��U��`�=؇+���_}�����C����?��w8}�-�C�@+�,p���9��=Γ�:���p���{�����{�'�cݐՑ������B�Υ��*���t\�a�c�XO$զ��>8��z�{?~7�翸��^Į7N`�Ӄ�x�����m�7�jK\/�cA��ת>l�}KUXMVR���t2�S�(��:Q�o��hˑa4�^�%K��"@�u$�*�϶��ʂJFT�p�V��:ҋ�����߯ڀ�<���mP�J�}�6v�6���
�=�����]tP��.B�6�9PY��a9��E:!?���;@W�ވ�������y1���?處�v~�.�a/��7���P�ˁ�-�_,��+��o§dǖ�˴��J��ql}�[�~�����	w}�[����smPG��A�(km���*t5�����]jf.�s
�WR���"4�9X���V�J��aH�-Fk�0������~��'��J�q�>��ݬ: ���\�֎>���+�V���M�����ł�?A�
OBlt*"��~�HI�������k�_7���=�N�t=c̶wA��u����e��ij#��@��ն�i� b��y|�0����s;Lm=�07 �-����G�`x�����Ll�`����Tw�!>/^�i۹ρ�t^�s;;`�VJ�u�*��W�lJ�o t�T6U*=���K�M -%6%>_C�9�j*�qK����kcDKQْ���0����y�k+X��lI|Y�Y�bDs�afgŰdXh�ޜh5QU��]$KjK'SX��P�m�s�Ά{�+B3�\����HmX���ĵ�õ0� ��M�/VݍW?�o|�>�r�}����}_Y~0���qn l����W�æ,
��ap-E:<�����.Bw"3}~�����*!J����Dh��2�z�(7�G��>ju	ՙ30�7k�p���������s�$fo�Nǋf3��|d��Gf�𘡪�r����d5�U�'��$>`|��?���%L���1��!>��w	�w	�w���U2�o��R�}:�/�RW ���\�=����こ��3��`�kN�8�j����L<O�NG��tt�ƳT��Ntr_|�<3\Z����G���_�?�o}�&F֎����aN0K����M��?���s |�-@���PN�h��$/Q���~�/�� g�,p���l̍BUg�>����������[��%�IODdU���&~0�y�OKĲ-p��Gx��������7�ī�ፗ_��o�����bۦ�h_Ԍ���H�ID\VB�����PTgaa�2��P��XЮ�:�Z��vo�ѣ�UO��?{��W.����|�8������q6<�f����jnj�96�
4�4( �8�W�hJ�R��������T2j�]�iLT��n+ �v�Oi�)�iz�%b����*C��Tځj3���ÅX�}�r�I ��j+H�Q!�QɆz	���d,Z�f	������&���!owDE#>.B�*�LA�T�д���s��ݜ�^pY�r�@T2�2/m=%$�)�e�ɒ�q�%H��� 5���t
$�溩΅��LWGM;Pgx�=��9/Uו���_��\Hځ
�5 ��R�社�tV$�� �z����!��sLe]y>� ��<	\�ȋ��Ҋ��7 4:"�zӹ{<~�"��PC�|��U�ѫp��A,]9����>9��O	EX��hX<���HȊGNy6�[���ׅ�c+�u�6?}�����ￃ���?��'|��Ǹ}��߽���c��Vl�u[�f~3���Z ��<,XT��Rxv³=O�[[.�3a���9��ì!j�@���iZG��D��^'Uac0S���E��Dh,�H�&Mo����*Uoۓ`�ǂS�V����TB2����*�2�#H�W\���E:!����~�w�����A� 4�&��� U5@r��sM�`^��h(Օ���
��׫�n݆Z���,�ڎO����y�J�2/�r�d�N�S���k|���A�Tc%6ey�/��%�(Q�A�~J��&"�� �G��Z�]�h�@���;	�m�*� ���U���Pi�)�I�OS�@��Oy^�)�k�����&�n�k�����3�n����X��z��^�G���Wb)��#,��\��	,�c���!s���*�*���Ve=��5@�}3@�Jn7���e��O�<^^ɲ���"caJ��+���8�n���U���1:��6a�ݍ�ra5�؉�/��������?��^��el?��k��/X:��o�X���&�60	��Ǧ|l�inz�
u@LM*Vwc�8������Ol�ؙ�8��"^����O?�{���~�G޽�o��n�s���|��w(t����'��˻҄��^N\˼t�*m0����(�GA� T�kz��e��%���C�<�����h?KM�ri�9�O~��1@[���N�TSA��cD?��j��=�{Tm@ǎ����k1|hݻFѱcM�{TP�N6m[���#����w�iw�j*��
D�W��V *��.�Ӌ��S�Nܠ�/�������1@7��9��t~�^���	�KD��UXL��0,
�W���
��T�ގ��_���ǻ���z/�CP�7L]fH�g���і��K8�+<���x�$�Ս���Ģ��eU��/���KL�D���f�siH��@`TBc	��4dr��E�)�C\j>���#>-�+x,{^@S{��h��:�����-|���>�X���W #-���� ���E�����hj�Ļ|�m���HH�@W�02��������CZv>��^!�����9�L�{�SP.�m�˼@8��Å�upP�m�8���+��1�u���W�c��O ۲�$ ��HDQc)��2������k	K��7G�h5:����T��J��P�e1���sK�>@�ʭ �ZP�W�-��VE��.��/ⴐ7����vd!�(� ׇqeh5��Fc[���Z��#�4a�0a�z3�6�0�1��lC���\�� ��!�c����� ��F����{�\��/@Xe�x3v����9�����kp���x����қO�8�
��yp*��iN L�C`Ah�)��cY,�I|�Eæ$��|��≈T����ȒjL�G`(�mvƨ7��&����|�i�:H5�A��r�f!Ow
g�B�,=��q��4��-�q|�N����4�2���f�5�O]<"n�X��+��3K�ai��MB�}�SH�[�S#|�|��S3c|" 5�v�zx�h�!U��)����<�{8�-�橭��o{8�*�/;�%\l�"㺳�:b���6��r�i"@{fb��,T<�n+#��T ����m~�c|�����:6�ـ��D��g���dL|j{�%@��o���/�Qa�K$c��H�g�� ���:>��F̃]j(l�a�Y��%�}��Q�ф�][�����_���_��㗰��ݧ�cぽ�u�F''�9Џ�'O���G�w�n\��k/���������؊���Q^Y���8�f� &-A,�;�� <�E���@���	�ʤh4����X�|X���8s��u�E\�p������ÿ��9��g�fow����߭�+ TJ�S�b��p1*�� *E�n�bI�}J�Oɪi"�a��ʔj�-�~K*�m%�)�~J�SЩ���TH;Pi#�n+�*�R�U�j�.0
H%�à� U�W�I[�Tu����u\�H����^j{�N;���T��J�R���4��$��,w�Ӵ��귂TF`��������
�n���o�<�����/��� Y��S�4�5�#"�E�����<O��C��S:�d>5Q9��Yh����U�[���*���ᖪ��T��1Htσ�������%��M���1�45�\�9������K|��x����ƻ��µsذyK�t��>�h"����#&=
���H.ཤ"�ud�`��5�sh�^9�����O>��#|����ӏ>Ļￅ���N�Gz{z��c���]Ձġz��"r��=��^��|xt���Ԛۆt�m͂5!j޸�)0�O�,BsV��>Kl�K��8��Ũ�'>�a����n6'�,��d<�����'���'@�nJ�N�����.K�X��vB4߻ �M��%�����Y��a.0�	Ĭ� �,�=M~	P�4ߩN��ږ���l�-.A�D=J�jP���/�`��1�`�vP�"����R��� �G3��$CZ)Uo�çd?�V��dE���"i�9�JB��P,#65 �C!�Y��5Up��T�մՌ	Z75K��g����_���V�UˈO�J�S�*��J�Tz���X8��RW *m@�Up����T�\���ii�׮�� @+t.9�J� t�յXye-�Ы�%�et����T��v�mR�S����oUp���+���㻴�g�����+ex>eyo�1�GY�����w�b��5�xa[/�þ�{p��8�����)��ŧx�����w���	��Z��u}���D͚n����p�u�-=�
�6`�����Xy/.}������?��������o��W�!�|��p��9�]ώc۫G���~L�߁�6�)��9��RGoi�)����=IGC��SӶS����`9O���zE���;G�smr>�yA��á�C�������"ڪ����C`�'5B�Ob��&��ۨ�K:��:3�.�W�ߞ�up| �	ģK���>l�N��k���*�mj���z4��D���) �*�Z�JU\����q����N���Tz�"@7<ܪ ���u�������f@�ځ���ХgWb� ]� ���d���`�����]E�K�+��b�'d� ��Rl�:[/��"@%J�Nܚ$@'�����ؕ,�5��2����b@��e�?���k���~���%K
�;S�Y0�=vs�`�h��T����^>��U+PY׆��b�D$���5��HM�GV^)R�s��0���H�I�ܘ�$ed��%ck&"%�Pw��}���,�-���g0�b��-�X��ck��;�ѥcX�j-��"!~!o�~�����!�Hћ����89{ '�7o����{y�q&����������~�م%��	@db*�뚑K@ǥfc�$�����?��=�;/�A�l�GbAP�z����aQ��.���_|�w�@�qw�OD0rj�P�\
�� 8/p�������)JGjеk�'x=\_���,��?t~	�×�Uh��S:z>���WVa�R �/�|��FN5�IW�V�Qm���
����z鄈 ��Z�h��-Gq�_�YT�"ⳐPU �(o�к�d��z�5с����2�`@�MF����oJpN���M�O3CE��!�fdM�{��е�	]G]�qwc��V>�0�6�e�|r�ڕ�� �;�.�����/��|���y����D�HlέK� �ش-�R��ϩ��}u<lJ���"���.�l����5�Cw�:M�l<�1M�(7��,B,��@df��"}�tdΚ�=T�q1e��aBu��;����	nZ��]��O�>2��+�zx�x�JoX�-B�-N���x��}���T|h6���?#T�E�����9�6�sc|� �L�����Ȉ�s�!�����)>�c��	�/��=i�ic���&x��ylo��s�q���{�v��>]���j����4�A߳T�m7�E��M����6�33E6�77���ӏ��w�����P�
�v���~n�i�1Mu>�ȑaWd�?Lϓ��R�
�t�&McAlza���f$,
�a��x��Cx:���������<�_|����s<��=�{�.��xW^�����s�_�&���
����_|���/ ��˸j������׮��^��{p��q�9rN���.�8��;xX�����ME|J$bR#���o���3*&� MBAB$
P�����g���}=mؼe=�}�.�í�p���#���Lo�~����'��jgwG8�ħtB$ �27���)��@]�TD�qF(JCi{(����,S�7	>i�(ؑ*��M��금�k:'�K5\�d�E2�t>�B�:9��A$S���x�EIgEܗdM�/�I���ē�����*ˤ��� ,X�I�TG{�����+ u����͝sܯf��*�������ę?��p+�O�KxJh;�Ju]���G��n<6��]��<>�9����������� �ω�d7��\y.d_�xL>D��[�����hڀj�/���~�@5�Z��H�Z2�j,P���	�����{N��=�Ϝ96��2'@MP{�D�tB���Ɯ��������~���g�zo���<{����cϾ�X�����㑔� �k;,>1iQ�ˌCr~
��rP][���.��\��;7c��8�n=��{��s�/s�����O0���~Np%��3��TD�� ����K�4���Rx��µ%
��p�mCf3,aڐ
��F2��	Lޗke(�87&����eY�kJ�qKLZ�MT���T��2�D�tL4�M3�Tם���8�l��:f�M�|��	� �� ��X8o�{�qYtb�ܒ�ڕ?���'@�߹�2�ў0�a��1S��*��,��5I[���,D/����b��7�xU��k1xhc,k��<tl	�X���ߋƝ��h'D�=h;jvw�V:#����&�L�O�S��+ZC�rZN�V��g)�XD`��U[�UTȰ*
�|J�T�)�Nh_K���N��huJ��dAk��M\��� �NnS����u�X�̈ ��Ԁ*���� v�Q�]]��Dz��
F�i�Y��
���b���2:�˪"��,s�Rm��z�0�Si�G��e�~9F	�e޸t<�2���U���vI�S�yd��X$�/�Gp* �"�O��z�}�Wj�	=-X%�xL�<�~Bm���,8@T�ay~ko�c}���jl�O�\Y����"F�?8��d���S�������^Ǎ<��ｄ[��*�~��||W��"^���x���ƻ�����Oq�����]��#���.��?��s_���ҫ�ۧ���Q�x�(v�u�^;�5/��r�hɵ5X|uB���.���"��a9U�y��$R����b��y,Ne(�}V���d�vL����+��%��N��:T&���o���풌4��X�/�x����X�2� �k��{V����-(���z1����[;U\�ʣ���FCۖ~��� �G��f���B����9̲�>@��{4�6�t�Ţ����Ӆᯇa��Fյ^�"�@������Vl~�9��b^G1����7�b��I,>K��RW|��ZL2V˔]M���0����0I\N����X�oO�c��:�t������V^D��Nb=?����b-/��7�	�q,'>�]��1�v	���1D�>2��b^ܫn�Q��Q��xe/������=#7}��o9��ݬ�����ΈJKD����t����j|�¢J,L���Px���M.Q�I�$4ӑ�����B�">1!���FFn>b����V��e������w���]����*��`htZ;�PVQ���.<{�Mlٲ�s籀����dde���1Ý�gdKP[ۄ�$�R�u���_�_��'�ظi%�J��I9�sn�BR�p������ Fe;ݽ��&YO>vt���/v:��~�{���gW/X�v��\/̙�T@r�*Q�ӈ��P8:c�|�Xπ��ꗷ�w�&/l��wa�	,%<�\��9Hp��U2��|N�?�TA�k�&��6��K+����e�dM�%�� ��d�����HDN]$
k	O�x
�%�Ɠ�,�!Xx�,(�@!�Y,�N�ċyc/፼�7�BiZ�"�����U� �Y�%��L�M�1��Y��F0b���&FĦ	q� J�Tք��1,�,`J\�8������f���6��pw�s�;�"�ښ��0�`!3�-x��c|������е�~�!�W��t�����>|f|��kb1�6��a���A�B�Dt�Ǡ�)=e�h�pG���m��j��zF��t��#�� ���f2)FӐl0��Ӑ�7�3Qg0�|��`�J�'�nۙ���Kģ�"m2�&�ߵ1���������;{޲�������q���t|`:��߲�ŷ��o�O��\�]������<�����@jH��#�;N�>���������쎙	^������	���_v��Q{�$�W�����.�Mfb��t�0��8%D;e���M�1ha�r��k\�0�����6Z�ub���`�<�Y��':g��A���6%ǟ�d�0���R�z���4���Ԙ��(5$�ϟu�d6�b������?��)�&"�HR���o�����
����_�]�"����Ǳ���-�ţW��.�eL5��˯~�7����~�	�z�7����|a�6�X?�5ˇ���7��
� )1�񡈎'����B0��"������ ?>�Q!(��B}^6j�r�T[�M�V���p��M\�vΝƃ�w��W�l�f�s��y�"��Iϭą���0�;+X�&&���"�<�C|��^<b.��_�UUl�PA��S��T%z4��J���"67����cr�Vp$�@%;*��`Hzj���Q )���M�,�d7�������Â/96هd�h*�G\ɱ�X�2���_�c�me^@�ٗ�=g&1)@��>�Q�E�P-J�i�l��(k�aJ����j3�r�y-�X���x�2�s*�E��\�y�΄$#*�HfS�מ��t|������̳��W���:�*��30���ުݪ�u�2;~���-aaaGG{����W4*RڗZ#)!gN�ǯ��>���?�w����:^!o_��cG�clb-�(,MCjFB�	���BLJ$��c����̢LT4V�1�b��Uذk#�:��7��ƃ���.�?��ƎCېU��w�$���(�[2�=P ߥ��C�D#B�V!��A}%��)���|�`.K�g]
̚�`�m�:�a��u��T�������D]��}ˠ� m��g"L�ST�[U��4Z�
�E\��_��YI�mOT���I��h�W1�%�Ō�X�j�V�E�4�N}�� I�&R���ItE@[.�<�����	�}�&�ݽ����6��� �-
VCN��Ǻ���(
�ku"��r�U���d��xe
WԠn]+F�<p|%����
����I�n&47��nsA�A�u�����R-�U�]ٺ��Di�)@,&�d*cvJ�A�J�6+���X��Vr{�����mJ�}A��vۆnB��~�� T�/-��e��Ҫ��j����о��������e_қ������c_WN4ףi_ώ`9�H�����B��z�7���,g8Rmͽ-�,��n���� �9²�����Zoa%�/fY����^��[�j�M�_���~z	�.����;5�p2z�o��Hu�s�/��ڎdď`J��T�h�93����Ֆ%��6��!C4��n�a9�:~6����9��š����'��ħ'p��S8���蜚|�4�||��9��o���a�4�� �?ݍ�G[����������q5�����H�4�ȍ	�ܜP�%�,�f����2i'����s!(��(�� .	o��+�_�R�y\ʴ� U3����SB���\������g��.ϷT��.W(�1��c�2i�K���RUp���`���N�>�� ݀UG7b�1tnF��E([ـ��,��#Z��C�Dg'�y]�,(���\$ï�Vmgt��߇���� ��L0^݀5��a���ύ�]���M@�9��������W��|�XwU���k���)@%�/ |JUܝO�)��,-C`^�� �v5���콜�PW,,�����!3�e�u�}fZz>"#��^���	BHh,�����HMM'h*��چ܂|��F�*�G@(I�M�Gva=�6l���0�z�Hpv�����=}��o"b�����_�W���j[�`�ؘ$df�#$8����(,(Cy�뚑������]�s�{/:�Q�Њ��z$�"2%a	Y�O/A`x<}����s<��XΆ�k���v��?a�B��T5��ҍG�ޏ�	;���� t.��sT�Є��V���a91�z�b��.̽m�8��{����5vs���3����2�|HVTй�_ri���c%F�Y�H����Oi�/uܵ ]�@�QB�J�C���(U%<*�Y%@��z�&���,n�W�̯�Q m(ANE�� :�d���>�) 5$>�%`L�L�FUǝm�9&ħ9LPc���V^�1�w�9��n�N�C��]� j��D_ԭ���'���ǯ����h��+�cO��e�Ľ=� M�5ߛuu��%`NM��uA(l�B`� ��@�g��<+,(�x���-�3Pk�C\��pC��Xh4I�:H��D2љ�?e\���g0ˍfb3�y��w�g㱄�)��㙥!޶!>��	����8��8Z�cs|do��	�O�-��>��5��~�R_X����Y��������s�'&\���s��O|=�c��s�=�Y�Vfx�d��p���y��8�Z�ĸ�4�у|]�Nc40�Y�ϝ�����As�[�zz�&|����W���]Ė/�/+��σϩQ��'í����K|��V��*
�^Q�"`@xږ�£:9�]�ߵ'�����}����5���?�������g8q�Fw�B�`%"R�]	��a��١����<�<w��K��w������*A�ҽ�x��gxt���م�˖b������ft�W��8Y��H�CBl���AP�Ty�����$�(�ߗ�h����h(�Ae^J�T;P�'q��"���'?�?��+�_=7�ԝS��D�=�4�
N�Q�h��D�a1�P���;�8t缠Q�G�a�<D	�԰ ��H0*���&;箪�
�P$YO��I		���R�bKډ
 �f�,�%�tJ6U�A^O2�Z�ʶ�Kulj{ɰ:+�	>e?Z4�����j��2/�(!ǧ�nQ@%����Oړj� �}o��tB��i*S�T˕yy�w�y��s� 
*��ʹ��ud*di/+�0�h�)�D����NUǕ�Ծ�|�nT��
DU'Hn��`U@,`���� �ESڬ��a�<���׌ ���A�����nh�?���a��.�ו�܁_~�=|����[����}������o����b��^T�:��IFH��H�� "!�DhbV"�y��/Euk�wax�b��0�����蹣
���\V�8w�,�w`~�?��֐NdanG:�൸�+k5ր��
�ó=nmY��/�<��[4�Ü 5kN��E9���R5kLV��U����Y%�rcT�EZ�
<	Я; "<�7 ��H�2�@��J��֯%��~��~�#<��=�zpi�U0IX c��Jà[�Y��-��q^0\��Ҟ���b$���,�A�U��6���e�~Wڷ�`����:�P�-�i�@��E��"��u
�G�u��PV~Pm�M��f^�j{�F��Ԭ_�2��� U�)��V����zP頨js�ZG�����<@���l����qNc��'� -]_��h9Ёa"s�t�s� eI�X��fؕ!�����������{U�~bq1��Ò=����2��������},�\<2/�X����=S�D��t�q�t@�CT��j�REW2��f�e�)p�cA���@���r��0��D���K,�9|e���x�*˓WY�"ϱ�x�e�|�i���Xuo����Í��d;�?ކ�����rw=˲�X�p&l�$�3����c%�[G��x�0z���Q*'_��TV�g�3�U��,���! �qQ����S��U�q=-.���̿Afϯ@��4�!��M �%@�y>�y�P��+�J�R���va�٭Xul#V^��=+�h�0�&;P����}�l�c$*��{:�@� C�t���^,�?��uX}���8����V��\{z)6�[�-�'��򸪂�������#W`)�)�\qu;^�s}-ʖW���;�k�m=Y��g� /�]#�H��AJj6#G�3&6�a��H@ *��P46.�ϥ`!��W���W��������GJf�ـ��T��L@G�>sQ��j���(��FMcaW���R�Mݾs7>����}���8x����@���Gqq.^���5Dh)�ӳ������RԷ����ə�H�*Drv1�Rr���@pL�§�gB"3��Q����:�@A������u�EG�J��##��!	pp�BTL:��W �����Fu;���3r�	P��3@���b��I�8�Wy�:�CF�xH�-����_/g.�n��Z^��ת��T��5��A~��U+�7��D��
@�ڂ��e��8+���'o�P�xH�-l�S��#^�Qߝ���8��0ҁ.Q�� �gd}���!����>��OS�C�a�Ė)�i�d
c3�{Xa��-l�����doDU�0����  ��IDAT?цډV8��b��5��:q��\�wO�D}��RMש2���*��И����9ձj|�9%��+�U�?椲��T?��Fc4%���h��E%V��Zf2%���כ�4"-�Ȍ#<cd��I��6��J�IO��t0��j:��ᆋ-�;�ౝ^�5�k�����!>f|��9��%��]O�`�#~���v�/���+_W���-�ckD�����,\~A�~���� B-�PK>O���~�����_x��5;��Lu:d�{s�qk�-�������q%A=�X�ϳ�T�Lf��t:��f��Lm�n��!z̍�ga�^|+�������-x��G��S�@G�Ò�7�`!����!V8�����N��g�+ӳ�aX��h�f��>�	��Qw���~��ϟ����?�W�{	�6�¯0��`���G�aV�L�=�T���+��I
�L�����G�[��/=z	�Ξ��+�q���>�{֭�hG;��������h--DM^&�b����PD�b~�Ė;�厤�@�gơ0=y	�ȋ�@EF2Zˋ��('`���������x��������3�X��v�ce� ��6n|�`K���[>g.�	���S��z�ReT��S2�%m�Qk�q�A-��=-6e�OyNz^u#��Gi*�h�����KP)�������J�G��j' �fC����8Y_s��.,�K���A�L�rYG���X�Iޏ�O�� �`�P.�}G:>�����!�X����ڬdHݧ2�ڌ�� R��}/�\�/�ZD�2��999ٗ X�#�E�jk+��z�X�T�%���\i�"F�Rɂ�L(1��3����<w�%Vmmg��\�a�d@����@�l�`e1ɉ�x��-�������W��~����g����-��p��NL�^���
d�'!*��/ZР(?"4��!�Y���TV�,hKOubx�0&6M`���8v�N^>E�^���q��%l>�)�YpN�C@cB���ޝ��t8�dý/��ZV���
x���)pn˄kw;s�Е�9�raA�Z�f��=V-�|�S����bzy8��;?���Y�w�7&@�I�%@�ƋR�W*! ��@|J��;�tD�_�$w,h�ĕO��'��S���-�~�r�����k\�h�?����X���\$�#y
�E+�Ǳ:ԬkA��A���Gǎ4njC��V�φ�D�Y�Yк�)Z��]U��j���+P$�$�
�|B��QH���RW(�JO��T`(��O2����=���K���&*S���^r�v/R���,��D�y�:
������1�X�	����Z*Q����rв��
���`���ट��F����0N����z@G�!rH2�,��^ǲ��**��,��Y�b�ew�ʲ����q�[��)��B�y���C,�K�OzyU�$�$�� El)�J�R��]�{�y���!G���҆�����K�Q1�_��k�I�d"��<7�0r��D�6˟�;c�ES�Z���i�;�Ƌj��&�����uƍ��J�BkB'�I�u���yg���>�E%�)�|.��@��3a������ˈ>��˫4ð�]�ޫ������PU��oB{Ξh7���)�2���K�s^�s]g����N�^������vl���/H5\��_X��]�U�z�%�ͪ]߆�=�;���뺁��&�� @��N.�ۍѽ}�{��*:��s���@��%�dB���̋{å1"v��X��k��+ ]rq%Ʈ�f��������6��Z����l�Nz��n�2�v�����j�X�QTY�����
���_�B��xy���>B����4�Ӹ~>::;�d�R�� <&M���7���<����=�(,��]��n�>/� T@��EOD��GsGJ	���j#.>M���\�?�@��X"8(��eMM��QUY��{��Ԇ�B�&� �� �)DXl2"�Θ�X��ȅ��H������j6	����6���BQy;b�����.lD\r!,m=aa�y^�wX
�vs�0�����hc3���5 �Յ������F�+ά��5�$�\^��+�#�/t�N�b��/��S3��`H�s�MT�*E�J�C���d@5�o�:n��A�>�lhZ�R�@T��,�"B%��ZM�[h#�P-�z�\?��9lA}��%q0������L��Г,�7 t����g��P_B�%>��>�Q �5�	d�b�����~��� �P'x�~9�HjLC���n����@�xY���\�/��O�~�+wOcdm/b��Wך8̩��}]��Ժ"
V��*
�l�g6 ���B�5�!�Lmq�sb���j;CTXLG��tT�뢜�@WY3��?	��4�H��,��OG.!Zi0M�v�$Bk�ҽV�8gg�{.s����ڙ�M��ن�������e6�t���s$>����}�/~⅟���\����.�K=>���fK���\��\������؛�k=<!X��4U��)�=���b7񹆸%���#���3�C;��L|���|, �$@;͌�in�EP#d�����R,[�� G�υuV0�rY����KC�t�@�dh��`��È��N��'��*-��),l��ۿ����~��׎ ��v)^0����ٰH���@��Ec~["�P�Ƃ�Ww|Y��,KFf.���|�1>��s|�����f�vlڈ�;w`�����ZX���lt��1;Ui)(MN@vt8RB� ���톐��'�XP�Y��LZ,Ң���"�&?m�h��TЋW����;x�W������Ǵr����(�z"~Dȼ�N*�l/mm�΀����2���|b��[e@I!A� M��S�C�'D�1x
oAj�ꔈ�H*�.*Y;m�O�)�FGF)8
�$�*��f?e�-��sy�T?�	���Y�yYW��ud��ab4���|
�w�\Py^�:F���v2��d�
�|=�Qѩ:tq��G�	o�H�}���z��Tu\4e�i-|%S�`g;�9�<�6������*�F�+���ɹK��Sh��:����汼��2�#�5-�? �4��
.��${�9�c̶����1���l���#\�Xi;����V	���;��՗_�ˏ����+�q���݆%��PYQ���\��"5#!��o�"|�P'�a���2�4���R�wԣ��	=#=X�n%��߆C��؅�8s�,��]?��o�sb qޘ[���Y�Ӝ��m�p�͆Sw�R��
1���KG&�R����ܞ|x�an	���g��~kޘ��4X��ä�h�����j�(z��k���۬A�q�ڝ����@��3� :� ��hZCLJO�e��I�W}ν�2����p��Wq����$q���kPA������N^7��hG.�{���U�Ծ"� ���Y�eyhWڶv��h�B��u[>뷴����Z�j�i�)��ț(E.�(�7Q�i�I4
@5�o�����>P�d?�2� T��7& �TϕǂX�ʶR�W����� ��d^�q���dI�U���~��3�Њ�����v�^^��;k1J-��B�e�Je@��~�g��{���㘸�I��}t�,��L/�!�����\zY�L��*����s�:%d�B*���]@��Q	���Ur%;�s�e<���s-��c`�-��=h��!�d���l%B������X�D�D˩>>G��=�h��Q�IG�����]%T��}�d���b.�ЍQ^_�!.����/F��!=��,�Ju�+|_�U&H�|�|v��*Kֳ�4�x�_��ˣ�d+a�v��I-���b��k!.�l�;п=7j�o(וj���T�B�L��RWޛdi�='U'D=�5 �D��E7]ލ��U�� ��>���:T�mA���gI�6H�м��� *�@�vwadw��N�	�H����o*=���͏_�	� T���dP^�/��'�� �����i�{�@��&�TF���&�_���	��Aȩ,FCW;j����W���4���a�|4�΀���
�����a��r�������U���nh����~�.U4!*!a����V-�߲�����>�6��ޏ�&��܂�*� v٨(�Fo//��-;�o�AlX�/\���q��9l߱��X�����<�koZNbS��K|�x�3"� >�)�ǩ�K B	Β�N��fd�H9�6�1I��$Ly�.a������|�c��T��3VN^H��ǣC��QwP��癨�����������������Y-h�Z�R���lˎd[���؉�رcgro���=y����N��j9��{g��ַ�>����:���!��
�Ѱu���9\|п;��mc��q�t��~o-��K�.���t�}���#�즴��,�L��� Tò�!�j�?$hZA���Uh]���$B�De�dA	Pn�N���t8T��+�Z��2�� YlAu{�\�UT�T�D� j`bC���1L���	�I�ijNY�[����~���>�	.q�Ng�(�oHEFw.��Ѳу��4���.�3�W�᏾����x����|b��)&2�kb6y�K84���E:"J�]M<��D�-�U�p*��wV�k��Q���x_4�١����zh��%@uQotUƆ(16@����H37F��ҍt�Gp��t[��XcD���,�Pc�tw�[����>���]��}7���-~��=l�SoG����p�o��k���B��\,T���	~����)Ì�f�gs����1���ܭ�ugS|�@���~���d�����1~��:Xb,��b��s,��[�b�� ��0�w�� ����}��Ö�Ĩ9�l�PO�9����������uA8lk�`Z�fu���V ��_�@+bX���Aa8� ��0�V���I<����k��wx���c��0����R�� X��.
�, ��!h,���̃�d>����3�ߙ�2��ՠ|f�����,���}|�;�Ƴ�?����^���X�|wFj�0Z]���rt��%;MY�JMBAL$2#B���@o�x!:�)	��(JCKu!j��P�����Z��M���Q�;sݸ�:~���~����*���~��_���QI`�����A^��<\��.�E5m@�,aο'7"H: ���S�Oow�p�Iɸ	�p���~>�$M�P7A��R�$h�I&�	S�U~^�Y�J�Q��FB��׬i�)�{�H� K�����
���O�=T����r��9A����*��8e[r��y	9�j�#��-8H�'�4�,���zr�z_�����X�� R�)�d[�O�9�k���	�ʭ��r����[��:�RXVۑk*mF��\�Z˶��q��h����1��BP-���p$�,���kFX����z��!i���`ssi[o�0�����r����@�Ї��=��7냨(ɐ���
��pw�����d<p8�w�/�M��hD�)��.%
�9�(�)Fm[-��B��ǰ���c����p��������u<|�!|��}�	XD�ٚ���tU��e���p+�C_6|�K�ގX��T%<FJ�:Xסx�W�u���y��+�]�{sa����yW��i0�HSPC>��3T/�FD��nk6���b����h�tF��z�=� m� Դ9A4�#�_���[x� }��۪�An"ð4j2��T�8�%�p%@cF*�N���T2�Pz�	���89���,؟G7�����m'�T�G�ܞ%�F���P1�V⯖XlVl֣t�e�u(ߨS=P��d.�ꭀQ ��V�2�A�T˕���	����5@�T�L�g$�Uy�Z�JTz�1C�R%W�~T�j��ޫ��,+�hA��~�W�ѷ�T睂O�}���: b�h�e��70�2��9E�H��Y��g�Yq�I��	H@7q�Yb��eU�Vځj���QI�l�l����@�!|9�תJ.��͈��)n[ ����ni2�RU�A
�F���y�`�qK�?��A"���$�d^�\6�>bo�)��&��F��6ѡ��T��3|��l�0�E��cLA��G0Mx�t����u���9���|�PK���N�x�2���kiK)���<y�s�1ŘF?��B��\_�)^9ON����*�����]W�|*�r�Ni�Y �W�ɇ�	�y�t^��n]��c����	�\\��#h�Dê��� �9�2��W'@�d�?���Q,\�����o�"8��w���4���y�~�,��g\���{�~�8��F�� )z����c�'�Y@�p,77��U�2񹌍�Oވ�N����������ܧ���UP�	w� <�^\S!�\��فX`H�2�@t�9��78o���KX��T�=��)����y�HjH���>�}�� x���5�]e@�G��|t�c��nB�����֪6�		HN�QYѐ�X��6���Yٹ���AVn*j�15?���]�,�bh�0Ǝ��g	�,�ajqK{����������#���kj,�Ͻ�.z���N��������?� �����������]���j_y%�H��CMc�5���	Զ"4>ξ1��B`T6���N`blzu��
OW�Ϭ������;ZeE�]C�`��,�}��B�&���/4qŘ�����<����
�W�8��%�c����	�p'޼���v1��d?�}���V�ՂS��s�MP����.�Z���?PY���O.b�?�
��9��@�@6����L%25mA�S�$�{�A]/�=����eH��
���=�\�����<L�t�������1�*���џUW��z�j�I|�ۨ6�.,�8Ǻ�y�7'��H��FF_>���}b)�E�!T	Х�;x�w��o����.��_v B� ��VEæ>v�I�ڭ�~Z�ո�.)pmLմ�M�=����|�/S�Q���� 4:��^�h��Gϻ�Ȑ5"B��gb�S� �4�G��H�h��!��|=A��?�].�di��]m���+> 4?"8���kɀ��a��%N�〿�����%~Nt�B��`��1~�d�_���5���~�dI|��n��&�U$��c��:��ANx��Mu���X�9,I�����l,p������y|���M%0�seAw��_����6�($����^S���t�f���$
����3������	�>�S��Ð��	�N�"�jq����ȏ�����G������N�t���ݙ���
x��k$�C�Ɇ�p�Y�Ȇ�L��
�3V���ȶR��������?������o�o}��x�Wq��s�Dou5�k0�Є�*t��#'M�J�Gat��C��oDx�"��	A���T���5c��S,�?z�<�~?��_�W�_�����_r��*���W��g���|���#a���D"D:"
��RUp���
�V�{�*�^��H"`2��� ɒ�+0j`��S�T5�� J@$�� 1T�Re)�:��,�d?��!MP�#�����=U���Q�ON$��\2}	�*0�3��dX�c!���'h�}H�PP&��H�:��|��d�����x�m�����tj:R�����:fcpP ��9�3&&J���̡�'$ĩ�A���"�(�@��ܿ&ii�*�,��k�˼@S���F�K/�����q˼lK�-禰�k*�k)�LIJV��k*���gcy��A��g�C���H��/�OH�<��� �������R��6�26���9���\~�Mtah�]=������^��&H��C�,GBJ����h:��0�������K�S�p�+��hD�P'�f�1�:�ͽ-��v��+7�(�>���Ͽ���_V Չu����g�-��]&K�4VǑ���dߟ��r�-7#x�ޓ�-��`1{�aו�����(�ÐT�-PPi*�1���aK���l0W�CuB4��*������3S�yH2��lH�\�t�������nO
�;�`ޚ�CEApoH��/��/�����w?�<�2�f�������T�e���H��WDý5�w�pR	Ѽ�:�-��r�]��1q��8;�v��ko�g�U{O�zJ���s2&��)�~����:Q}���iRQN����	�nT˪���f��گ��~�W�TCMvT��J�\y�A�T�m��Pm�R`Z��	U���	N%:t߄B� T�˶4�x��\��T�BmW�U'D-���se@SS�U�+��GV���QE��'�w48!�枖rӆ�F+��
@���"E�)˥��T�yhF-��6�Gn�p[�-� t�ţX多�ki�) �6�R�Tz�=|{GM�UQU{ȧ:�IMY~ ��	���S��M��Z.�}D�L���a���xrN�,Ӣu��aT����/�|*�c�Qp� ZG��Qi��� �x���(|��|t������h�ÂO�)1������(���P�=���G���~�Sу1�!)�էf~ǪJ.����="�8/ml��5c�<:Tڀ�x���.��+Tt��S�y�,�й��;����!4o��y�GuB�̀J�~�S�a�8� :z��$J�����C��:����kG����r\e;O�sg>��<�=�>U���Ƴ;ؔ!X�C�Ml?��-���o�7�ʂ��G��T��6���)�I��+2˦&���&�@����d,�����W�ݵ�q��������xՓU0��Sm@]���ũ;�cC��ӎ#;�Gm}�Bfbb&ff���5���F"?����n}C;���T��>��R�������*����*Z�2��A�T���}['����G��q�>u���������������/x����O��'o�{��~����|���&�]���������td�����:T�5"���e�h��ǩ�`k�
���T��h92*��iT|>"��n���p���q��/"����0��s0�R�� o�h��E!08Ee-�)n���M���/c��9���?-�a.�qԃoV����S����)�v+��!c;-�(�է*����'��K� tE *�@!�����%�{����zѸZ���T��ć}�}�h���L�tg��!����S ڕ����%���p���lj:
U/�zċ��YUp�	�;Up`jkK+X{��2�va�p�r�s�<3X�"N���֓���b���b�����h��@>���>|���x����x�� ���d�Ş�'<�R�Ғ�@�֜F�&*�:���(߳���E~ �S<�������G�6�^��7@������ج%@+��F6Q�cd�B���a4s]�ۀ�)&�fFX4:�U����*����9��t��=�}_���	?�qď	ҿ"B�m��a�-���<m�3k�̝Sw{�;��^N���~�����/}��5?g�����:�u_{<bo��V�8�}��`�\˖z},Y�0�q���22��{� 1�'B�!:�������͖ƨ�5C��%by,Qq~p�arCT�2��X����N�t���Sɨ�ġ�H�=$ -��u]2��Py���u?��ZaXL��xæ!}�ZYtʄ�x�ǲ	OB��6���Lh�1��{ݾ&qex���w��_�������_�
��O��������~��o�Ʊ#G0�܌��Ж��f����MIBi\r#B���� �x#���^.�tB*�E9	Dh6��3Q�����2��7�k|���5�ŵ�.�_|��a�������yL���caz�D~nZ
�i��bo�x�����PPi*cr��"؏`��@N2t6� MU�%�4p�U�F;M�ۄ;(xi�����2/JA�d<������ �-UZJ�£�&%s*Ǔ�����,d�:���O: <
BU&����K($�W�ՠS3D�� P�rP���� PB�AJH���D��S �^�D�^b�C��R�V[�X�����T�M -p�J�1}"[�eRY��&[�������4߇�'�E�/���&�	��Dޫ��!��)I�]Ʃy�#��'R32Ґ����S��)�2ll�,7��f��2���\���Mx�#� u�h�FCK	r���ODZѝ�H421a	��)<άDd�d��pk�j��׊��>̭�c����=��珫N��=|�<� ����p��:̣�`���^;R��؏���19�;"�e�����XoS�'D�+�6Po�L:&��,:3aѕ��|�T2��vM�It��y ݇��|������~�	P݃ �!:9��H�qS��o[.��e|�w�������w@M҂@��6* 5���{{��9݀̉ZdOՠ�H3��ۉ�Q��Gx�A�IM�[���Y��@��6�S��l;?���Df3*�*�|�sz��g5����*YM�TJ�SBڃ
%*�PMȼ Q�)�CU�t��ɀ�v�j���3�oi*T��}tj�)ռ��V��֣v���ک���i�T����bH�2�욦�'�o.�L��rՎ��d9Y>�g_��%��d?e*�%c���|� 4%�����V����,���%�)�@����
��)C� d�o��$�|b}�t��2��zw��T���2����$��A"uX2�R]�H{n�S1��#O/q=b�1��{��j�J�*tJ5[n��||� ��y�о���P,ᩍ{��Tb��H�%s���E����tB���S�q[c��,��r��"�� �>����1Z��e�@�
� ���(Z��K�Ώ�N�$�weC���?���Ut��46:��o��+���.v�8����dC�ѷ�p�MMܣ�е��ԘL��s�it�\.Upwn��#���ǎ���{�����x�nc�]~I��j2��9�1���a	�����8��)<���񹟿��#�0����ʀzGx�#ԋPUp�֖�;2���.U�6:&��/(���?\\}� ODe�����ާ ����h>|c�@�aX�X �O��2��(�Wð�Vw��n坨o���`c�z��=�Ǟ|�xۻ����@UU5***��ٍ+���ܹ�(/�@Nv.��|`ldoN��S������bd����]�c8}�NAPL�3K���Be� �{gQRՅ��L��*��EM*�)O�S����x4�aI���@n~5&g7��U��V�zc����ZF��&T:!�EXi6#>o���3'����0�h|I: �4@���!9�#���0,�/�^{eGat�y�t/A:#R�q~�?4��{�@����^͇g����,�DcO�	�f��ج9��R�6�i�b!��#����4��aՒ�:!2��U ��*���0�3���l�$�;؆;�>�n)�
�1DbrG&�'�P:_���!]��KN t�,���ٽU�����o�/����Q䰐X���BE��L���*�r*�O��s�v�|��H{Q��N0����.�A��*
Gif *"\P�I������M�QK�U����
��F�("BK	�
c]T3L�aa�AsM'>�FSD������(����q�����]'K|��o���;A�n�;��{�'!���po�<�W����'A��Et(�6&ߋ�WX�|����b���ys�����6�U^�+c�ٚb��[0��4�9n��1C��c��
�C<�!#����];�����&�M��c��PWx�x�*�&a0*��>*�'î��'�Y��S�$�9HZ�E���1��y�]_��d���h���>���<��ê/փ��J�#�B���@�>���d3�0��I�5�P��k/=������׾�'o>��{/�z��-ܼq+��km�t{�Bh{~�Y��|���aHT�L�WUo#�P�?������LGB�󁿧=��=��1Ahi����+t�=H������"������
�>�8r�?3=�	���Gtz��� ���
�[����{n��o���0��S�!v�8��l�=-��2/�����BQ�݆|N2zI��,��eii(��Cqa�ss����2���Q֗��63*۔� M�(���m�T�'��������	�������8{���ʞ��S��	#�� ��H{Hi3)�C� �MB���%LJWڤ�>5X�6�S0�1i�.�LMue9f9������<Num	d�>�99>y_z��Ϛs����������/h��D�d>��p4�, ��\G�����$''��p�:�gT:&�����������������|���{8��3����p$���>*��8^�}�F0bӉ��dg���U-�h�nB�H7����������k�\�ӷo��C��|lM�ɏ�CI���6^��bX��Ú�&��B8��#�p�*F�j���#a���Up�΃�p����5]C�f��=]�^B���lIV�O��t�P)P��h ڟ��� =�Y �#@%t�R5��ct'*�jO�AC,#��|�U|�˿�~�m����h]�TUp-��U\�DPC鰭2
�mH�i@�b+�ь�J.6��(��� ���h����
���r�-2�К�l
4%Jl
<U��S�K�TeR�U���D�hH������^S��@��E���b@��g�3�NɂJϹ�T�) ���T�� ���I=�ZS�r�]��0E�-�2� *��Lhw8�2��[�U{���m*dNGsOi:��t+Upf=5mAY��T��J�[i����,�/<���vU&t��X|vS܎�[�9�}�T`�zE�D�2�J�C.��K�������1A�"ƞ^�8C��� ��yHS�U֑���v;#�ϰd����c�I��1������x}�վ������`H���G�ڭ�����?<�c�Q��j�CR�@<Om��RMW������2Y� <�! pJ�sH���
B5����uԼ��= :�����ċg@���\TùM��w@����@�f7��Ϳők�׵)�_Ǡ����2����b��eMt�e����q#:O�}R��$�P��w܍gwUT���&�nn`��:C���'>���8�;!����׎A�������Տ�,����^R?Х[�6�_�� ��&����g���X�O�'���`�`v¼��Ҧ�����5�[e8#��: ��jPW�� '����kDfV�XP���Dlb<����d敢��_��Z�g��Y����`f�vN\��"��gy.�G02>���<��x�w��+�`uuUM����btt���x�g������it��`p|}�*�[\���&��FvI�c������T����{��Ω��6���w	������TGd�6�ə�
��_pB␘����4���7��X>u]�H�σjd'=�����3���)�=����'5 }������twH�S�b�|�?h/o�*���@���P�����4�{/��~M�*><�����DUW�ꐨVz�m�`!�#M����4��,mKB9�59(�MG!���I�ÿ��o;=����P����6v��w�}�3c����	3����4��`Q2[�ʥ4�F�v\��`�DL;�w��9|��_����#���*��ט���L���é9.�ipo&d�܃S��L8���]1J�ZI�0)�I��s������E	^�qF��9J�tQc��j}T��&�(&@����� �&z]�we�*F��:��~+CLؚ`���	�U�PWǉ���5C<�����%^p��K.�x��oy:�=�O�~��{8�MGk��h�7]�p��
OZ���%4w��MBw�T�����cm�m;+l�[b��Gx<3D��a��&�Gx�#O�y@�����Qon�r���^�sFH�7\R|`I�G@�4�D��@��[�?�JI���Qj<P�8�{��B��U��viG�ał�EwB�k�PBl��~$��,���y*N�ٰN��t>���:Z��"���e�\N�&
�ޖ���"<����7?�����S8�s����ճ�pvgG�F1�ۃ��FtUT�9?�i�(M�Cnt8�ÂO?��"&�����.B�⁔� ^/D�y#&�Dh�7l�M`��k�0��308#C]B$�]mH�>,�U�[{Ks������.D�+�[7��͙x�ri*Up�̸��3}�U'D�T$0��� G����H�& $�k�A.Hi������lO ������L���Z\I6R;���S֕L��S�`�;	���e�:���B*8�>e{rL�@ٟ��/�e*��>%�}O��t�8+')�)|�Y�4��8":~D�a���`*�D����[2��}y- ��u��d��,n����\{�Z��T�I�?'��lC�/�T�Uf��P\i�)�M�f�!�T��'\BZޓhRB<��SB}�z���<?PX3l�����g7g�y�������pp�z�f��3����\���� >����; gĤ�9I*ZTS���;�pG�ǰ���͓�8yi��Ͼ�z�:�N�1ށЊ�d+����n�����8�Ip��o�~� ��p�p�-C���D�l��׫�!3u�_h��`��E *�pͺ�`Dt
>�Z�l�Pm'D���Yf<����Ym@�dD����G zH *�����ۑ��8���]����x�_�+}	O��,O��is2L	g�Ȁ �+��sK:�&k�A����1m���(]iF�ސh��1tH����To��Y�ٓ6��h�c��T��h�!T�hC9�&Qy��M�PѬ^WkA�1�!K���R�)�c������,��6� �@Q��|Vnԣb�N-�V���e{R�V�+�tjڍj������&ח��v$d��S��+m@ei�v�3O.`�e���>]w�	�F�iO/�v���y��7�<�Mt�mMi�څr^����W�6�|���Q��$�Q�?�Nɂ
D�J�,�Ή��z��5�s]A��!�=�j�#����~f��0�c�{��}z�[�t�h]�yH�I"�PӶ�<XmU��6Fd�?O"������4��d�k�O��dEU��OsOr�OI��UM�~#�#=�JO��T!��,�j�'��&��<�S
�<~���>>�xmd*(�f@P�Z���\w�f;��%\|�>У7�c�c(����8ڶ�� t�~n�~� �,/���>Be�����)Э�[|
��8� z\ J|�x�N�}ZeB���Ob��q�t�i���ul2�x�m�g>���g��8�I2�'n���+GU'D���t@�i��E�Tý;��#��[X%<5ñl`��6��	\}�
�*�a�e�2��a������e�X9��cgN���Y�ň�J��w0<��TO�2��G��hLl�������B r�[����"��d�,(d棸�? ��(,�@bF-R��;��ݓױ�q=��>~�_}�������O��;C����Μ9���~ǎS���7|�;��ŋ�F0=u�����h��Cm�zPPU���8��! :i��X���:B��ai���D$��!��EEQEz��<{v.��v�BDL
�xM�fWx^9���2�{�:燑ٔ��@��B����-���l={�/�Śd@�
�m~G/�w�YUp?Sm�ϭ׎�q@U�Oi�y�05�����cs�ԇ��j���b �C9��� 0SPE|ʸ��h��#U�z+C�HT0����C[ Zڝ�R.�*�2���.���q@��?��^peP�y��1�E�x��o�2�����ve#k�eu
��;��^k�G~(������x�k��o��/~�6��ݚ���l��&����MvoɀGS:��3������LP�D���%�0,�~��&��Mq��3�b�Q�
;�;�{��E��ʈ�R"�D!�E��裐��'�N	�2������N^�1k#�5ú�1vL��GX#�����r�q����	�˦��JD�Ǹ���:Q{�p�H�^���{���e[��!l�p�co���q+3��V8bn��r���xLcM�O�~~O}fF�17">�PGP�[����e��`;G��#���^0��~q8�J��P�Jb9%@ˢp�<��1@���SC̚Sa���Q���C��Ra�£�@*��Ra5�Lh��a"S�#�m&�������#%p)b���)�l>\�_�x_�t����
~����gq� }��}x��#�q�*�=���	Luw���u���L�������"2�R���
�B����@	4� x�0B��B_g������#�s{;3x�;  ��.������35ԃ��)�	'����j��p���Ԋ�$2,�amΩ���Ց���.��Y��V�EV��J��*���TW�j�4�(�
�J�,���R�׌ͩ�����^��mr]��`K@%���T�:;��2������bOU�մ��ITګ
"�Z��v��39f�5d ����T�)X��,�����|��/�������CTL�B�����_�!���T��G�(�/`��ӌ�ɂJV�+����L	���\�Sb�W^i�*�'�@�!��dr�
��O~VzPДj���I�g��^��\�����B���U/������L�����Ξ�8:�QzQ&B]�`��{��v��u0���1�1Fp�;b�ÈfD%�{�6�	���|2�3���T���5m5h�k��䀪��}z�����}��<��C8s�j�����t5$��h!���j�p�)e��r"�D��<]� t��G6_���J�ý�@���,T u�o��p1,��TDz��Г긝i0�sˀ�2��T�2�4ν'@��Z�B���@u�8����
��:�`�J���9�^~o��x�����^�Sע:�-)0����@���Ҟ�h�3i���fL�l��`��z4���u�/M��ؔ���-��=�8ً��^4JT2��Q��y�e�|�sz��	��m�a�0
%;9Ȃ�dC��Dm{���|�k�)� ) �{�� V ��ު6�M�j����&��v+�k��Jh3�������֣�|�*'m��r�g T���5��){�T�*��K�AD����`U[���{���kmGDԱ��5�|2$�)�o%۩�����ΰ,\_2y�%�lG����f>��"��d/��� �M��S���?M�N�8ƹ�QnW֓����QB3��~�GN���6Cz0�j^���S�f&6@~2	6�	ehz��,� ����-��T�O�&�����O��[W�Y �;Uޗ��!YMi�)�OA��T��q&���~���u�б���7��ʛ�g���,]��ԅeО�ch�D���;Up�`���:rO��_��__���q,�7��[�Xy���o����
Ɇ�Rq�����1��:B\J�>��c�O��Ǳ��.����~|J��-��[�id����Sb� @�x�����@: ����K�q@�=�.�H쾠��VzP]x^O��<+U/ ���?B��{D2����8]%H�_��_���?�������1�^Q|@��;���=<��3{h��BzN>�ӳ���x��f�A�BVb"���4d� '��Df}S7���QPZ���BD'e#!�����ElZ)J�{00��gƩ����)�N����?�������?�3�@���)��������c��'���+W����=�:��|��W/������ʺz����~��v�Fxbj���]XO�X8���?$�IE�mhlr1�C�0���������g8��WX���<ػ��?2� ?@��X=s���h�%����m�ptm��̫װK|�|�'@7� �?_�w�?ҏ��q�O��Ё����`s���~�s]�"��7��<>���T�$@�׫P0��B>(+��P9����4��ҳmE;��u)Z�ץ��T�U�Et��]�e�|x��d��;��(mɁ���fPB��ܐ5����I�H���Ԙ�4Q!5�k��$l��3c+C�;����Nan�$�9(	GhMb�ґN|�T�d�U+-�81���.xEB7�����[�[����y����8w��&�R�{b�M�������)p#B=۲�K��r�]������x�G�%!0*$��aP��7X'9�7ѝ߽7�c=��w8��RŦ�(#�	O�z["S�����	��S"?
���@�!L�x��,Ͱ`e�u;�
�D��~�ؘ(5�����>�	F��3�:8M���6N�C8�흱1�I�g��[�M�o��b���&�72���.�����wX����|/��>N���n~�m��jy~%���q2C��5�B�Og�%{�2�f9�0)�à_	��(�1�K�3\�n��X���'@aNh�LW���<�O�����9{͇�i,�f�v<֣�c�^
�#���T�͂�X�F�a���H�ρ�\�ʀ:�$§:/|�M����=�8.]���݇D�3�����V~*�P]����4&E#;.)��Fd���n���u���3��!�*����b��!�H�	���qhW{��
�D9Ã�n|Ϛ��vz��D&�`ED����dr��l	k���\�vj��9ב���bec��vD�����`�m�É�p�a�F̸��/D������ى�9���g%��g���;����km�k;�+رݟ��٩�e{NܯLe�..�j��)���Z��� ���p'�5��L0��e=�g=�����:���m�q�)��}��:��z�T��::��+Ydn����2��$+��ϻr�nܞ?�ho�^{�~d�r�kWnߛ�#&��������p���3��low.��qJ�����;�x��!���H��R��ۛ�����+�_O7N�q�y������x��}��1)�dmg��6D��{k�8���m9�٨p湻��	PgB�Nn�*���}$�������\e#+/�i��AXlA�F�<����>ËP�P���:�vcvy�gvp��	\~���^x�1��zy�𪈃k[\���m�'�a�p 6%���`C|�MKu�b�͕�q� �S�$Dj�=Q��A��>��+��`��2^�weC���v��#�!m2%+I���}�0ʁ�p��*�P��i�9�ɀ��j��	>��U�D�O���>>2<�	��Sۚ�� ���7������k�[�yv(̫��?��$��XU;�(�ud"n���,(#{�����n�v7�/�@}q
mh�ހ����!L����=�yN�*n�~�*"N[�V�l����r*�;�j��ۚ�$S�wi� �����h+��1�(��D%�P/�a�F=�%�)Y��.#:�I��+p�rҹ����z�=����6Pٷ Sڏ
h5����6�Z�#�����,'����q��}�Eb�e�)���X�����D
��ϮR�xd��4Q:-x#L��OI�넧f�OA�d@e��� T��j:*C��,/�|N��?+�r}���IX�},�*��HuQfok����k{Xeq��� �p�G�3\o���g����ב�%��;ɞN���.�%��J/�M�Q��'$Ӻ�bD@�2�<�T�}�!m6g�����BeU�v��k+��N�|*S���<��gL�8��ٶ�AxjC�9@�
�e���)����)c�����jB�zB�+� ��:����C�-��K�P^Oٗdhe����~��'����{�2.�~]3�{X���j:*���y���n�Ȝ��}������$D9&6%�����0F��)"u��)��&�^�����y󸦺-�)�Ʉ��� �y�86�g���U1��6��x� =F�JD���xch��.��yl��n�"l����+����h��u켸I�nc�M�OM'D��vȕ���>��{� �@FP*���c��5�H6�y�����<���h^i�y(<�6p�t�W�7<�}����I,�Am{����������%� � ��JBTh<"S�����<�Gf"9���uHͬB|J	�YDt�q7�����{	�՝HɮDe �G��=���K8{�1�l��Ͻ�[���o����W�O���������_zo����6N��xdy��\%J���O>�k܏'�~
|�Un�WV"���2�KO?r�*� '� �����7���*�}����ڃ��� $2� -Adl>�S����b4֎�p�	Ctz��rzmS]H�͂S�t���Ꮙ�8������Ϋ{�Q,ݖ��˘�����ZlJu[���S�]�3�T���~+�|N?!�����T :|�� �D�h:r�RQz�H6��R����,iKEas2
	�">������,!�2�ׂOy]��ۦ�Q"Up��*mA��04�n��O#XN2�S�Ɣ(|����� �nh�1����q(Bkc�r|_RG��?W���V4���ko��[�W�C!,d�0,�V�&���Ļ_|	W�C~G>�RYH�M�GS<Z��ژ��87�0,�pkφCc*��{������%e\H��C�ȏ��q��3=��?B9<��a����@��!�͉P�jk� �M�P)UUy�E�b���<�C�1;�lsN9/ˤ
o��)�--1da�yK����].;MX\���U[K\�1�Ukc�!.[ᴝ1�؛���)�ؚ⬭9Nۚ���ذ6�
�_�6ł�)��M0J����H]Dm7����3e���tZ������L��
>����}%��":�Kp�K�;������C~Fe�0���^eU��aЩ%@%"T53c�d�uˎTx�p��Wi�ٕ��,Xf�l4fcY�|����υ�� S�	{��L������A��Rx̗�]�a�,�O/��Bq��K�-�	o�󶪲������Y]]ř�m�,�op�]m,�T"/;ى�ȈAb�"�<�� �ӟS_?7x��Ĩo�B�łzTx|���4zU���@��1<y�{5�ċ�T�$$�e)�MK+�ӆSb���\�=����KS�X�Ô�5�af�ud���Rp"x��>��$��C�Ѯ���~�+b�q���q|j<.�SBp���3�9��{�Yַ!ش篖�#l���Ö��v��������5g��I��ך�.���:�D{��Y�u�l���he'���k+��[��^�)S���ٷ:&��b��WN^Cs^_����V��,�a�l{W�=��4���d�<y<P';����\uKB�I�1���Dqa>���qxi场�z�7���a��@Zf�2QN��4���� ���~l�����Ӹ��E|�W�譇��[�F�K{��bMU�)�NO�Sp�)�-Æ���k��B.+��l	�*�P	��r�}���Bg��O���U�{�
�3�p�k��b���������g�A��5����K�']!T��B=BR�S������\��T�14��P��T�`�7G�@O�2/	@���������S��Ͼ���{x�K��v��9!0#@M%�ْ���Dè2�ϧt�OU#c�^��&B��UGD�}�H��@�)ⓡ�z��c�h"B%d��m?3�:�Z�Ӽ?�f�OT�}DVnH�R�������/H��P���g� �5����P.��(�r�l���4H��ۮ%�ж�ݚ�^7�O��㔦�]���=���P����\uh$p�&����~���"��_?��W���m��gMs�i��!��2���Z2x�SYgB��`Y}��X���3�궂O-B�_;���\���w:&~P�kD� �q���*S�}�s�n����/찬�N��7��*+*�F����k�T{Qm�]��T��*���� �!�c���e���N�Z�,!C�H�F�_���u%�
� U3�1�c�j��yٞ����o��'�>+d=9�O�,�T�=�_�b"x��y�{�SB��~"WP�j�����C�}eG�O�{�����,�&�7Hx�yH�9���Y�8���XF�9��(�;���oL�6�Z�^x��=}+7�c���IT�_D��I4���q@�Ύ)����������D���q]������1zu����I�l�����;�z��~;�OTuF��I��Ox��`����xGo%@��uS�߮��Q[�bU��'�΋+�Jl2����n��x����3��2�XX�#�>1�p�jc)1��\�E^E�SR���ȸ$x�"8Dz�Fld*2������,���#,2�фZ|b���Chl.<�Xp�����{�0�B��[܈*�����s;�~��g7p����ٯ����]���������W|��W���h>��d@�axtLuX��)�>�ԓ��A"�����O�
�}�mԵ����C��X\���h��GHt
l��`n��BaJ�zE��?^����!<����[$��%!-�
���ȯ�E�H?ﭣgq 	��p��P ��M����p��Yl�xۼw��������0���@������%�ƌ�S�O��t�Q�8\@�f5
&��7��b�KX�/�1�=y�i(jI�7@��R�6�,�˲��$��aXИ� �o�}3�\ځ~PM�� 5> Ps.������BHE����Н���dOW���kmh��Aϩ1Ԯ�#���' ��0f�~�=���������͋(�,�Kv ���Z�
7"T�uɰ���6��0���M}���`E��	���q���aB��y�0Os�m
�⎄x7�E8!���R%�BO!��D��A�K�VI����^��\�\7� ��zEƺ�0�C��Hv���5��2�2Q�eg�cvf�c��7��y3�t0�q[c��5�i{s������y������$�c����F�'aIpJV���Ixv��4cp�=\�AD7�5<�bK�:�!����tA`�;\�\`���l4/���0*	�� S Z!���~��T 5iL�UG:�s�,�/�Pg�ÿޣ.�ʀ�DΝ�f��V�Y�͆�����ra��8��S�H8���B�/���Z��r��µ:�����>^~�%��l����8�����)�s�]������P]Y�<i����0�G "����%@�� Ox��Iw{�d������bd�&�0'�pe�ߖߡ��Q@�z�^�� `}W�@O"�]�E j!�OBF�SPBC�!! 3%<���4!��	Ì�tp9&S����&L�ٻC�{W�˔�;�-��j_w����0�1�9�� L$,�c�
��Y�9�����<�O���,�P��YnC���9���"�HfR���`}+����Vff�*�d�m�Q�l�f�02�Wa¿UsS�Lֱ��e;Ʀ�021��n��MԵ���}�d��i�h[W{�9ɽc+�� O����������CyOZ�K��~^���Bm]%n<� ~���{�f�=y���G *)
��q�)�DY]	��j��߂��v�.Oane'�ű�;�����ۏ����]G��;��Å�t�)Tm>�P��q�v����}["�a�n�h9�����"x�W h���p&.%�'*�G����ú�f���@,�K`>T#>�T;ОU�ax�=�%m69�!�$�PC"TeE�T>����@4k=�7$�Qn��P�$J�|W2ے�S.C��`���<���|O~�6���EWL��jS"��iT>��y����d-���(\���Z:�Xؽ���ӣw ������Z�6%9m=��GZC�	"�Q��@�(l�����
ɀ6�P����';�gd���Ɠ�Gվd'!�x�C!��xj75 m!2:	N���}�<�	��+�M%S�����|�Pyo�uG��v���#�}�46���	9�}@�3r�\c^����Gb��i��W1%<�^xZ��j�) �ж�o7$KI\
>���8��O��ǉC��N�х�UFt�YM����=�,:�$��|���*�S����0���@<	@5HԀQP�$���o��K;X~�����^K�=��j�
��M"H�8�ʴ!�մ+%�>��ن���د"{W(D��d?gU��w�SZ��%�$Y�q�s��E��d��*�#��,��eh��h�A���fT�W�lN��da?��-�̫�0,Rw푓X�� eY�2���%��*�Jt�>��:���&	O�= �e�8��5�wK�M@g��UިXye���+����z��S� @_V ���[ǰ��~�ۛkؐ6�<9O!>��Y��bn��S�M�����s����3�{��J�a�o�hwx���=�!)Q�� d��5�
G`dK�|�J��8�"*,I��H(@
���ظ$��"��	��H˩Ava#��602�E.�}`���X����.�od	�Nݏ��M;s���������w��׿�m���;���å�W�����ɛOcu}�E�������B���$N�?��^����O���P�Ҋ��"t�N`t�0V	��Sg1:����\PkG_>��`���b4�i,d���5^ޱ'@��Lz�m����=����}|�;���ND���.�z��%�8��%�,v_>���?,/o��Wfo�������&��!m�S�O	�n���W�д]���䎰0<��B>@�R�ך�����i(lMAZH�IfT���"BT����TQ��f>�k�`�Gx��}��	 5!̴ ����[�'�ӃP���Xĵ�!�?�S
����(_iA�F'zό�e�A5�0gA>5�W��k?�*��/���xg�n�f�
�-���] �ژ� �© Ԧ:�D�MM,O˚x�W���8���A~ t��B?��{C���D�a����a��o"44�qѮHrD&�%��y��(&.�LuQO��ʼ��t�3��5Q��VH�Iv�XB�j$�r���Z��.� �:�k6��a}�0ֹ�e�C8b��e�o͜˹����Q;��K��!F?��@�,Զ�-<�fsC�2��ݵI��Ѣ� ��ħ.��"d�����&�}�����
�tWe�i���D{Q�J�`, -�n9�Y!�O�dB2Ν�s���ЗW��e� v,��gÙ�tˁAi=�+�L�d?��GN]Xhu�,�#?�Jt��v�Ϭ���|!|W*���,�FO��n����n<� �7�q��Gp�˘���`��0=ҍ���T䠴0�)�HK�@|t"B}�����/�ѝS;�ӂ���\,����(����ވ��TXX�gX9[���v޼o���?nӛ{g'�JK A�X	<�jE�J�K�WZ2$�eNl�I�Y��@��:̉����N�9|:�%�#!5٧�d,��%�u0,��3�����N�{}���<K�ww�y����&�Ps�Vr��
K.�gȶVܞ5�I�O��|�\�)�D�!U`]`�L:;��Ց�'ة�h�.�kR�ؑ�d,Oɖj3�R5�����R��]��YW��Jc{'{8�9��e���r\�n��k�d/�8[�������;�}�}�&�B���}cKCxs��P/�g�;Ѝ7�y��_��k�g���� Ħ�!&%�Y��)�BYC):��9؆��6L.�a�Ȅ���fW��2؈��R�5���#��AX����z;ÿa�;��a�v�	��o�N��g����]���1�ɀzΔ�g����p�g���[R
ǡbX����@1�K`9XS>�����p,&���&B;��#J�v������P�T�g�SeI�s>��P-F;�4�J�&�E`�ƞ�����x�/�m}�ya0���UOL�l5nN�~U*��(�f�5(���!����B��YLݿ����x��QH|
<�v��q���n�C!����� mQH86H��]*��ǂ�d>{/�����D-@���x���lK�'�D����}U����TU��K���A��un�N��g���OD�(�������h�nꏵ��t���ϝ��'���Qf�w�YA����HS�?��9,��=��A�,���7yc�������n��>D�H���[�TӕqD%�����W����&���)�ns�l(��긏,b��dK��b���X!B�^=��w.�̸��)�� Q3/UeR�PA�@������Og@%K)�p���8�Qy-���O *�Z,0$���L*\��J�t�t7<���$k��B-�N�}d��� !*�*砽NZH�=8�{`�ǳ�y����gt����s8y���W ���9�?v�y�.����ug�ѧ2�c�f1~?�s}#ק�@�4 �R�U�N �����gg@O�yJe@ן���cK8��*����*�)c�nb�5�K�C� ��~�*�ɋ��/a�Bb���&�xA�wt��q<��#��ރ��fA/���Np'������fL�A��8�#ba����"�V6��Հ���� � K��C*ᙖV���TTu��}��S�iD��"���.�������������uG�Nai�VNa~�$N_xG��02}?������EB���_����~�����+*��/}�����7Q@}��7�����~�+�����.�����r	��R�OL�w|y�(�k�s
�5�&B=b��g�H3Ξ�p�&J������_�����T8r����5u�q` �71��Hȕ 4/�đC�����������8��il��P�/����[�K ���2�ʢt6%�F�7��T2�3�ze�[�(��C�p:r����MGQ�Ӛ�"��]S�6��A|��RՖQ̇vA?��e��.��B�dҫ�4 �8N���� @U{��(�J�ZyX�+��9���A\S
R�s�1R����.���ՅZF��~��B�V/��a� ��l]?�o��k����/����Idԥ �>	���l΄kC��:q�^���ɰo�!ZR`S�Kbժ<�0.Q�O�A�ȟ��b_�3�
�a��	�t78���/��qH�pE��-2�M�k��R�C�1�A���	�{E��>*�����dN��J"����c41�=��c�����iƌ�I�r�4�8i��Q�+x2:�F��	�ij�&~M�g3��c�p��e��~j��Z"��� E����B\�=��]���k��I�;��qA�~^ �%k\���&�Q�/#>�Bq�<���8���n5W��ʀ�p>���`/�ʆs6�i�΀�h�&r��������J\Y0�궞�,� �d;bN���p)�7j�݀؝&d� Ut��;=>7��S�hl���f����	-��h�+Fcu>���PW����d�� =1�1�{�Cp�7���OO��y��x�$������ӊ��y<t�"����6v�04ׅ��l�ly���
�@@�|��PG�8H�S�o��T%t8����`��Q@"6v�-�mðrsPaNT�V����ejIpX�ګ�\�������!��;4��G�?5������)�}w��{�n�r><k.��g��w�߳& ?\f!�M>/�s=	;/�{�ޙ:��Ù��+�� ox���?<~���g�F�#26
!�!�'^wOi��(��&���n�s������0�s�jȘp�gfe��0�y����Djf�b"^Ga�d@�w;o���l���jO�����[��+-U�-�M��������?�s�]\�r��|�ͯ 9=F�M�B|r,R㐞��GY*�JQ�Z���&t�chZ:"����%L��i��uY�NBxOF��1)=U�I�9+ -���҅2M� �����,�������z���D�f��ֆ��z�r=�hPڂ�����/T��/��[��� S��c5Z �ތ�N�Rp� �핪�*۩�9Hl������VYR�� ���T��V���I�6�����:����������򯾇/��/���^E��$l
#aQ��ɀ��¤%F�D�:N��
�9�M� h�f7��,`����M���V�������y ����jY#��� z���d4��n��qM��W��wi�g��SR5V��]*3*QY_e<UU�--@+6�Qΐ�[O��>�>�V��5�� T��}n@M%�) ���tt$	2���{U������u��o�3`�%���`Wz�}�8���r�B��S�1I��?���_�����Y6�#ʖ�%��^�"�y���E���ڪ��PmϷZ�J���9� S�� S2�Z�
>�_:F\���R *�QA��Sڅ�z�P��L�-��+'TT0(�lj��2�� rI!s�9�)���T�Z[W^��E��iwW��d?ƛ&�)�?%ȟ����dJ�G �u��y���j�
��MM{Om�P��+��=MgE#T�K������&PU�X2���C3��/P�W��
@Wn��ԥ��A��$�W���م����*�J5�)�0�Y���Up�V�U�|��~n{��@����]���� Tڀ�p�@7eH�'W� T�D-@W��:�)��7@����Õ/܇_~�35����s�3|�}��po�W�cxi{W������18z�2���GXY;���f�xE��H��DRLR�J��[χg-�
�����u��Q���qbj�(z��3�c�FW��Ǜcv���0}x�������^x�U��/��}�淿�G��&����'�3|�?Ŀ����7�V���������������%R���
DaE%*�105��g/����9H�,D1]Z׉��:Eg��7��!p�!^�����ȄO@��c�J��!]�RP�ߋ3�܇�㇑P��4��#�$G�=����06��=��)����#���^\R �|n�W�}Z~0�C֑!V�𻔱@�3"��-�p��[�H: R�����ߪC�=��,>$��@�&(��|��8�LC�`�;�=�(�Cq�ga�GY^Г����T&�� 5�<�f(�) 5V��� 52���5|���O|6$#�#���ȝ�@�a�=��m>D��}
�m��+��^�5\S�ri_���导���m�������÷.>�٪��ᩲ�M�p"F��-(Aڒ�FAh"����9�oZ��P�����=T�Q�{C'��ٞ���w�7"���o�8 �-1�A�����Pm�G�ꡎѠ��&#���Nu�^���D_ך��������6���#0�	�n�����q�7F�������c������l+��ct�����E���h"<���zNk�P�}�X�#�Rلt��⢜��
�wX���X��N�����WD��z)�V��4�D�n�t<$=�F�|�),����a 6,�Y��¼'V�)p"<�F3U�O������fI�YPu�+��n��r�-U��p��p��,�İp��BL����!�xu�����B\a�3�T����T����6EI(�O@MY���Q����Xd�I1��	@h��(�!m�X��e�?��7ו�������x�S�pt��.�7'3����N��^!�	@`�<�\a�dMlJ�UM5K��)�'��,U�N2x�D�dO�8����ۅ�u&j5H���tX�}K/'�;���f��0u#����0#彻�ܛ��^���{mW�C�}w�ʱ�	!�|��˶��y�C�� �����%d^�m��!�O�jȶe�>����$��`�PSw8z�9���>p�_t��"��0"4<>��pp�5��PU�e�Ҭ�LTUW����yH#Bc���	
��a�� ;{[xz�#)%ť�hhn@kgJ��� MFי�-�["�ޛ�v�Vî��~�� x��U/B�ӝߏ�1����*�����7�|?r?���o�u�GD���ah��=䤨�~Yi.jjJP�T�ڀvw�g�s�>2���J���!�2A����z�\�T�}�T�-�ߴ�d?�	��RF�?�|8���\w��3%
�3e�$f��5�#:�r�<\ϩ*x0l
aI��p��
�Y�̅�X?*a>���e�����#��,&AI�J��h��S��������"iJ|��h�ӕ�m�۳��:�������ç��o~x'ڵ3��hX�cޙ�Pӆ4�ϧ$�MV!g�Y4m��Nt��"����i� ��&" T^B%3*0�@�h�L�`�yO��������yuBe@;Ж=@5�o�� T>+ې��C�-[�S!�IF����f�^�ʂ
D{�����'�)Uu�"�W�Y�ߋ�����x� m�9Toԡ��] ���uGYn�"@Wdԁ�V1- }��+�E�خ��U�	�����,��~������������\�����d8�]5���,��s%�)����YT�)ˤ:��-�,c��U�o�e;b� ���p���U�9yO��JO%�(
�SZ�
��
�d8ǟ:|=���]�A�J{Lٖ�6�P͐.Ҧ�`TK���q�w����w���N�}�ލO	YG��L�r�mi�w�kB^Mu`-@%�m��9�須�W��P�H z���p�;+�n>~����}[9;���[�D#�&�Oa���9��k�Om�I��h�Б+Ø�<���S�J�[i*P�P,�'1z��8��Ӫ\�h���Xn[�]&@%zL��QUw��������֓�	��z��b�_��+�ܼ��G�O^�{t�P�W�)C�|@�]R�yhC^V֬aY�t��g߻�Ǿ�$.�s�;�+
�[�+���߄ $g�oqg���YD��`a�(�����|H���#���H�+@jb1�9�H�BBB�����FBR1����[���[AU� �Z���=��y�6!�����`��%��z��K�ʷ��_��������|�?�;:���g��;�ѯ~���=��dc���/��?��|��D��\�������1Զ�Ǭ��ۘ]��9M#��a	YȫhF��"*��������'��c�>�)����BlJ>��r��x"vb}�|݋�)�'�ai��#����z[/����n�_���D�-��B���Ax�?!=t��hVMe��7�dJT�]���ڃj����LUϸ���:���j�@�3���"�ŜnB�+�'ZО�B>��{�	�,5-�c��!�yݙ��2��$Z���^Ç�#!I�����Đ5����j�$=�
B�P3�Ŝ��1�c��SCY�x"0�7���țdAl��S��6��<9��B���%{�333'�Ɨ^�׾�.>�ʫ8sii�	�/A`C��S�ْ��L�ԩ!΂��t8�`d[�k�j`KK�P��X�	5�6�
�`X�����g���R�|�fy�=��<��8w��:��a��	�	��C(78�"�� m��G��ڍ��JC42�F[U4��Xue=!)c��p����0�M1t1`��A~�\6�׾�׻]2�暪��&&�"B�L�������g�-�Q��,�3B��҃l���$w�����
�7������ WmdK���PPòpVD@���$��TE¸!v=�p)�4��)�e�v�1���4؍p:��\�ȸ���p�/��B�N���dx�K��2�,V |�I��H��@�V+��+��¢{_l�b`Z3~&^p)��WY|Kc^����$��#�,���(̏CqN�sP����H�Ą !*H!S�����D�\=��J�9Z!16C]�82��{��o~�[�<������a�mG?�C܈Pw"4AQ�u��9��6f�&:��c!+3���ħT�5s��3��C����n
�&E�ahzw�&��O��P�yr{����
���a*!ۿ+d[ƞ�0������
S.�T�&\����F��҆1�^X�� F�A���u-x�,PKԊ���s���l�aC|�2�:���p
�3��P?xG��ߙG�/��y�z�pc���	�	HIKQ��O�G"��i�HNMB!*��x�aa!���@	�Z�(�(Eqe)ғ���f�_ז����Vv���}� q=/7�51҅���|�6�������w�o~���ȑY8�=�{+&>)�H�LDQv*����XW���j4wգs���}h��B~gB����L_��w��/�G���
������Jt
@���*��s%��.��D�FsU�Rׅ�t��zɀ����'�#2�o)|�*������`ۓˮl����/��V��̃�3�4�i����$�$tړ�TǕ6���S:"RONV͕P %4�\��P?�*�Pơ�d�	�%j��l_�_����^��{x�w1~~�Rc$Fe@�%ښ��$P;B4r��u
��	���Xm���9~l�W��u~]�FTP�t
8���`T��
�P��d'����@��x��ZA��z;� �� ڤG]�SB��JFT>+�l�6�{]wZ�Ӥ����?�H��RW��j�zʼ6�)m@������1?e�z��kz��d@[���z�S�ŉ��`�s�}c����˻,?��6�S,�/`32%���YÊ���'�x�6p��m;
�k|�!�_�t��sU���T;$� t���l�d;%�[��2L��Rڄ�,���˩`R %�F������,��Y΃qS�dG5YP���~�S��� H9Ҵ��eW��t��w�����N�,��2��B�yw�k=ٮ�6����eZ���sќ��U��z�V����gV�T�!��k��C���܍E\��}����x�wZe@�mb��ڶ�P�҉���0���J/��W�(�y]2�S�|`V���1�sHt�� �.a큙{��R�N��=�&A��j���.��ZS��gw���:z� ������_����	"#�q�p�v�_r��C�XAK:���64���f$e���9U��JCxX2�C�����<�%������τ�_��1H�V��"5�
��j����G����ۮ�B
�"��f���71����g��{�cU�V�)�����~���y_�����q�����D]C#>�����J+ˡ�w���+)Q�մ����ݣ�ZZE]g�Rs	�D�f��cc[�l@H�,O��K�������\b���\?���蝙����a��Q���"��P+x�`��c��o�������IU�V�^�|���ś�?���<��
�_�}q{OK��#����aT�V#{<Y#Y��@&��e~W
��.��f��K�����y�����̎Td���H�� ��LF,���F�!!�:�P��l�J\#CΜ����Ь��W�p�eK�p�F�F���|8�-۽(�1�t�!�h�>�����*>��x��gp����LDV� �>�5Iw��:�P�eH�O4US�*���0-	�YI#�E�0.�aѕG|�:ž0 ���a��	�f� �M ��B���o�چ����� �D_AZ���(�)��X��4F'���h'J۸��׶Y�m����m�v^�^�3}�J�j:.��{�f7ߗu��5�����m
v��U�G%�t��m��t[}��#��
����L�Dp���<`��S�� ���D�NϽȟ�ǡ�`N���P����25_.C����Я�e[�s�2��>���^�?6��,$��a4��C2�s,�.�*|�����yb�o�A��h$>;��Ӊ��R~��0�c��dhu�ܡ���o�g{�;�Cm<�R�^��X��$"�&U�K�Ѽ(dgG� 3�I�H�BBL �"|�	�@wx����e�b��p�t7bj�+�x���Obl���������y� 'x�{ 0�Q)�O���5�lMB-�,P��ƶ���t�����d�$�(�4�L!��)<2��;��u�\�p܏ M@�������"�!����^���k�w����Pɘ��q/l�s��`j.�\�Uv��d[��!Q� �1l��Լ���B�k�/����gIx ����x�1%'��q���FLB���M�C"�)�$MOVUmӳ�QRR���*TTU �(����-�GbF
�	L+�R���[����NV��3��[:���u���y�	ή�V�*��o|ȧ�������O����Lʌ�1��B<��cˎGLj�SPUY���*�4W���彵(�30������.��Uf Lr���YM$�&���[-�^�߲T�%8��K�m;�o\��f�x�r�Ԑ,Pɀ�����=YL|��c��Q���ZD��*�J�P��jx�U����-��i�=�p/���:��Ԩ긦�0��Gh"tGP�>I�ϻᩍ�����?/Ph�?έཿ�&^���q��wX�Z�Ma�+�aљ3ɂ�$ì)� ���W:!�9;��V�d@;�)pJTB���Z�U��'@�wZ�6*�T%0;���*d^����U8풱E�Ei/*�;� ��~�m�ϲ���Zz/)h�dE��	�fCe=�X���L5ð�\��8�V9v��t7�Y�>��Y�z�<�����m�M$*�爱�}�J�ۥ�+X#
w_���.�y�e��j*��oe�|
@%���6��tH�rg^:&��P�SY�h�|r�#�18�ud*�~F��c`�G�}<)�P:���fU�@����F"�q{����4!��fD5����������-P�~�d@�}�����>�m�ҦT2�2����i�S/�Sð�>u��a��*:|f�;ê
���=3��+�}D,�9v?�D�L'����k#�O��̕e�{t� =��qUW��eѓo�������6�y���Է����h[jEdq$|�}�������"�$U]蚘@��$*��PPQ���x�����LAXH"B���T��� ����l$%#/�]=����AFD�ڑ�V���Ie
�2��opr���Η>��^B?�{���x�q�����_�5����~��ߪL�׾��nGW7R�2��م��yD�D�����dD'&":)	ye�Mu-�;��?5���*�G�3��ѐ8�Q�6�ΑEԴ�"������#�}��,��#-��@MG1�x����W�17��:>tS}ab�ܡR\}�a����8��%�����(�^�P��?7���B��
2%���Q��jzý7@�/�� ��A�H62�3�ѝ�@�ߝ���\w����A�����9�%Fs2/˲��WA(�e�eHگ�+�#bʔH2&���Ď�	5f���� 5&�\C\����$��#�� ��,�,ԣb���NG��"m@�O�gouKmH��G@n8������{�m����91���4��G��&.��
��'���J�[�Ӂش'>Uֳ>I�Ӯ^ �KbTz�5-��y��2�*�EA0���z���-�!@�aT��|/X�y��u���_��=TF41�I��H�0E��!2��Phe�rK#T��n�������M���6��n�����^�.~��˻�y�N�r2�	�zF�Z����4�'<��gAt�����j�hsDD�"<ɉ�v��i_�	�|7�@?�zE�*��Yx't��BT��I���6��"Y0�R���"��	��4X�&�p���d4�cp��R���-d�����2�O�~�q^t�F4h���̈́Imz>���~�?y%�0"�M�o��hX����!N��}�
�ܖ
���4&#��B4����D$��#�0yyq�H�@rJ0�燠H/����=��x�s�|���e�̂$������U�h�AA�4p���%��@���9�n����� �'�6.2��	L��aakF��ħ1!!�p#�� K���Hx��!�ݍ���BPww���0a�;�Wy�����].�;>�Rm��O�{���LpvW�r�:V��U����z�����]ͫ*�Ğ,s	�G�?�5���_D0B�"���(�R �E\R<1��D>S��$R3S�F|�g��;��������AQ*��F"$:\�3u��P�pM�,@-�,`ʰ����������e8x;���:�:8�4�/���:ۑ_��`WXx��9��i�>�IEpf���U��!���R��؆�O6!��ٰ+��-qeS]�̭��m,7,T"l�A���7_�9�m��ٕ�t�߷B(QjO�J'D�u"<]�N�Y�������ь��Jx�*�F�4���<b�;�=^�����!J�����\�Ӭ�p<�k���mV�v���-S�BM��C� ��MW�}J&�^�,�g�H�����0j��~a�.�᫿�1�𓯫6�=|nY��g@�*Up?�i��
n�J;��L(��\�U�o���S��6�d?%���e�޽ ������m�*���k%�)��k�W2���dE�/��u��EU�w	Pi��E�lW��c�
�]�� SB�_�W'D-İD;A, �#0e\л��˛vZ���tr��Y�>����2�|p�޿���vYFZR����skD�	�#��}��>��2�یu�Ru0tW@�c�j�C�ZѶ���K �l/��T��j�<�	�.
��*��2�˲��ԧC��RUGUm%c\�w�*������OnS1�YW��C��x�q�9 }\z��c���6*�T�ׄ�%�c;x��!�'S9g�y��H	OiG:�8��Ĩ�:���G�?��އ�^�����K�t��k]h��VUp��	��s���by��zHPt�@��}c�����'2�o���;�=lݒ(o��C*�R���o=��/����a�P�>p��D`z���W����~tN������?
=�HH�&���P.�?
~ޑ�MG�_"|�b����Z���{����-hDJF%�� �$a����UC����Ex������|���9��nC�]���8���g�PUq��_�/|�Gx��x���T�ܚ�:��ᝄ��l�&'#<.���ȯ�FYC3����N �Yx�K`4�1H̭@u���O`��%<�Ƈ���	|���C3H�)ETrsJP�Њ��uLn����	i��pIp�k�;�.�����<�K_�_��\~Qz&[��-�@<7M�Na��s ��^�y�?v���M�>�����������F��9��t>ӺҐIL�ve��K ���|b3Y=��l��ħL�uf�L?��b$W%��I_�X��S U�@�@M���؂x��f"��� Љ
�-6��	��������}���8�>�	���,����2>"B���s8s�0����`5&ؔ6�R�Sڃ�sR�V�a��?vu�ê&QnZ��hWD��,F�1�dA��wB*@�+�!j���\_xd��?���.MtDx��C���k�TWd�(JO������3]4���D��j�2
�������:sC�K�Z���!��vC	C����h`���h9aZ����#�� iN�Hp3F|�5bb�/x�z����S��J����2���_���+�,R�O��$�T[��Џ1��PC�����gӜD|���/�퉰�$�	P��X�'�fHP��4���� T:'q|��3��h��I|:M�ø3Qu����� �I��&6����K�eS,��aRӆx�4˾��4�6�.R%�Sw��S����$D�%!�2�y����߼/����8���pf���V~ְ��{�r����O���
��V�r3���l��5׵�0���%�}�6p���������!�lLP3X؛6w�#�9������Ś��a�F�2�Ƙ�`M2�wŽ�5�������g�A0�g$x�Ɯ~:�лB�t�3�b�'���T!������C:7���I�tD$ms�]`��D�T�v��d@���A�
�tJ� )τ�DP�|fHv�0�Ey���"B�PTT��ত����!�����W�/�Â�C��{8���愧��,	O�hXEx�(��t�+���k���L�c�#k}�Z�F��u����`8��1+�͍EDq�*�����|dL4�no����M�AI(���`ߒ Ӛ��PU0�[��7]���V$l�˵�Z(����^�� � u�-��S����U�r����l ��my�AsUH?>�ȥf����%[hDѥ9����v f|�Y����E�+�51�6_�����
�w����h8�|ޚf��0mM�Ye4�.�+��>��w��7?���#�-�R�+>W-��5kK�EK�=�9Q�������봴O[V�i��S[�V��=�Jo�
@�w *�m2/m>k�4ò���#�}W�TvS�!�����,���:n_���v:$C�H;P5�~�\YG��2A���6�#����m7l6����.��-���x�4.~��}��{�/nc��U�=Ct���
�d�ϰl�X~~��d:�l����Si��i��|H2��|_��
B��\O��j�{*�K�A�Q$�RW��"S *����(u0+�Ń��>�ɐ�5m(�1����2�2����v0>�/�d�i��q��O��?�q�{��ٮ�dcy]_V1� ��e��Q	^뻏_s����'�*�y%:$�?����<&���G$k��ʀ�|�"6�Ú�6F�-�#j���>������}��yO�`�a��i�i� t��(�"ɀ
@�.c���}�z����������*��,�P�Mu��&.�w��w�Ǵ���fg��M ���`�eǣ��K'��0!X�ڊ��$g�")=ѱ�����W�b��T���^���#+�
��EHI-Cw�������b��g L���4&A�����lD'����1|�Ïp��yL-Ϋ�nϞ����E\�|_��q��>O�9�����T�\鄨�����O�&#2>1�)H� �J+PT]���O�����Hd!
�)y�*kB^U;�smC����`q�"&�GMk?Jjې^P��"v���,�"����
�E���}����.�� νsۯ��2���۫�z~��Na��� ����P���xy�?~�a��{�� ʖ�P� 4�7)�HkOCVG�:��m��,�3��L�C0C�y�k���d���"�%֞f��fF�0��24�gT��&���D|Q"��s��B��-C�"3��l��t�{#�;vy5��Q<Z���=�|�2�����ᇯ��_|�ݿ�b�;�!D� �EŒ�2���)phH�SS��h�&�Z2`O|����,4�ٵqЯ�ġr�,z%��'�
`����*�&Ȉ �0!�l
Yh#X]=����lWb��	NH�E���C4��E�a)a^n��JsT��֚ꠞȯ7�<��P�6�C׭�ul4$R4Ѣ/S}4��F�\��Dh������(p�B���B���ʿO�f{�=��wV�C��:����~�?��=��A������Mi����F|Q.��
�ea
��D�[/��{к���M�Mw^I��O�� �O�����p~4��,P�o�s7�s��e�s����\��l�x�,�r�ģiU<,�`��ϐ�;��D7%C�&z,�5�A�!���𜭀�#�p���И wBկ1	��	H*GtV BS}��_��('�[ÚaFYÌaJ̛�[�9�MS_+����w5�9�V,�ښp�	&\��a�Gx�����^p B�#+}�Zi �`��i�J,F*�G���~l9]+r��'�V��V�����)�������C�������n�g8��X�zĳ>C���\�+�>^�1߽�?�����Y��<
��6���$��������굃q�全��A���+�c�jz� 
@��S��F\r��vJ�S�ғ��������U�6��c	�����Wו�V���(�x�^��������-O�_y2<K��]���x����*�ƞ�W�``o =��޴��{V����QO�My�$���u
��=�H�F�l3��"f�v-D���am��`����V�B�<f���D�v�W�PW"ӝ u]���b9��Z�`q��j�p�T�!Up�&��i�Z�/�#y�q�?܀��zM������\����<N��f0��Ep�,��
�=[Dn%,G
�SڂjC�)џP��+P�e?a�g�A>tao��+x�o���~�,����������̵�H�z/�f�W!���ҥ�����Û�4���~fHaS��J��eO�(�Ώ��u����N�ŧ�d-U\���̧d8��[hñ5_����N��8�mh:5�6�RW �ŧ�K�?i*�>~F:��g��N5��TU�=?t�}hב����!A�T�U=��"_���i��>Վ��k,s=��5bq���H(ޔ�t��r1�څ>����*ֈ�U��B��
>Y~�'������%�'\��V����s�T�ն�\�πjڂj�]b�M��jB ��t
<�������>HUv�V���P5���m?�)����
N5��E5��/�)���$dٽ�6�}��s��	>� �e����?�MA�&�eHMTPɀ~6@���5���x��^��� t��cY��Z��8�{/��շ$@/`�ɳX��vw0v~�GGѸуf���j:���	�YBy��L�C��}��h�|?���������.�y;oJ��&���IM�Ϸѷ�`��38��Vonb�;Z|�h|�N�|�R>Fx���3�عI��\îē�����X�
��J(��z�n����.,U�W^�T�|{�0�*�Z%D��(�)=�2�|�9�����@T���!J���^�����c8����2�.� �5�f�?�^�^H*N����>xm�H�)@aY~htBC��� ����`��1,-�@yE��c���rd�T#)�q	y�":BKl�f�":>>����6�˛0=��'�y��?���#X��������|�X�����{�)��?�#�	�����B�����xDD�!*.��MFt
�UX��r��4a|y����(�ER~��Z�Yގ��n�6!2�q�D4�O.�GQc/rk[�US���.t��ky�㍼n�pH�Fdu:�o���w��{<��׏c��֑�0k	����s��x��|�7;�8��"o~�<�?�裳����I}��q�ߗ?�÷ְ��Q�xn�{�"c�߻��sy-Yѡk�(>R���4��#�7��I�# �PM�IGrORzL�
BS�����r�٭�,<�`fm@���11�<jl�m�)�ԆLMex����M�]n�^��IC,a�Г���b�LV���t@�Mx����{��x`}禐=P���l���o<����M|��������dW��;��j��gm2ܪ��\�'�CU1����Rxw��5����h6l���h�WFÊ���x�V����2�W�uK�Dh�ϝ�/�D�f�}3��F�Bb����>���}����oD$y >���$\҃��a��CH��A��
-��4�'@uQE�W3j�&�(3�A����9�k�g��L]d8 ���N��r���$��#2�a�c�7,K	�2O�z���zeh�/�~������D �PSݲ@b����ꚨ���g���Q0-�aq�%ݓ�.⿛ѓJ���^U�M�U_2,��4،�6���|8.���2�̗��X��Dn�we�����lq X�5�gW����Am,�CBҀ���t�cq�1zM	@ej�N�e�}�~S,��é3�̈́sS��"�Y���8x�F�!�nEap��u�r�T��.���;�P�5�"mq(�
:Af�	��a4�I�;q=��P��LͶ����m��<��c�C����V6��J 3GB��0���	�(�!�	��_K;E��*H5&��͓��kCΛG�N��#�	w�ӁH��������.<N��Z����f�w��v�/��E{�p[<7�j�dA�[��M�in�?����8�C����{�6*Ƅ���C�,(Ռ�)�0	�Uf��6�q�gm�u-�cg
^'K{;�:9����6�0��pjj�k�&�aac�'�l��ޚמa�	S��
���3�c�klΰ�5��v���+�=���P_�D�?*A���I��oA�Rb��g�Q)шL�Bh|8��NPLB���k�"������E|&"-'Q	Q�����S^c=�%z"�5���oKGx_�;$ރr��C/��k�{�3l���Y��кD����"DOV"��K_oG�F2X�*g����b���ؕ3�ɠ&���4����uq0�ߒ�1¿A��h��kȿA������#��{�bff�T�bffffffFU��,uKjAwZ�j��t��|���1=��x7��7�}�|_|�s�%UWk������7�|1s�̕�+sf��[c�1ǋ�ׅ8�ӱ�jx<��*�"cB���D��D�|��X�"5v�g� >��{!�\/r/#��	��D�B�7[��w�D1�J�?U��2���{���.C�:�u���<�P1�Y	;B�Ig*�:R�ߞ�4��*	�fY0�Qs���Zo�N���0�)��lXRc`P��ˋ�������?�5~��?���-8煰���}WL�5�p�[Ra�>˩.����gL5 u�� Z��B�&�m`��"Z�m�F�DЬ��C�u�ݬB;�Y�qy�f�M��kQMh+�nD�j5�t�ƚ}B#��P�&c</�	�Ch;�OP�F�xWOu+5�8R's����LA~�����.�qPR�A��<��3<G�7ɸ+�Hz;/��p���˺�S���nB�V#j����CՉjO�q]#�O4k�� {�M����R᷻��uڹf+I�$���k�����8�a�=M�և{ئ=������B��ɴ��	l~��B�<�q�6�<!S`t��8-�H����>C(�"�Nr�@���d�O�H�G O�̎.�t�t�X7�}趕����P�V=w��{g���P3��*�.��-I��en7�4$S�<^F/aj��w��Ų��%uT5�)�m�Ǜ%H�P<�H��H�o���x.�<�	�L?3A�M�K��u���iPBN�9�	����,u�ב���B!�Qƨ��]*�eJΡ��vMh�H���p^�Jy�y=��^��r���x��]��=�[�A]��ݚP ��B<�o���W�\����1um�g&	�CjV��=:���j���[S*�v��e����$w���s����k��"��ߛ��.t�S6@�<e*����$��d��_�ǩO�a��9�?Y�����`�@Oh ��:O���f�6 ��� ���o(�@��)ਖ਼�C>k TyCe[��;O��{���V�p�~|7~r�z�c���8F�/�GS��ʮ̟��?1���Z�U!���q9����#Q�CAaJ˚��WC�:������,�������dBg&£�9&Aa	
M@FN9;�F4��������_b��9�8}o@�^����1t��g��5�������?���/�!���p�?1�I��(FBl:�	6�TJ��3�VTD��@qsz�'1����4���}4�@[�ZԄج*�fV ��	�UMH�jDJY�*�P=Ї��u��Z@�d#��^E�I>���V\�������X��!�~q��`�5��ޣ�|����X������B@G%�/Y��b���OJ\�C�Oi�N��h����{�xQ��R�\���4$S�})��"�v'S)�c���k�K ��F�3�0�* J�<�u"��j�a#^S��*�L4 *��&�K��A 5��hn#3#��-���<��$��#m���B	��dGsr��� ;�!������<7�Ķ4��`xo7�_��?y?��>y��6��G Hp�i0|xo<	���p'|�U'í&G��q��T���,�.�� ɀK���:���5���H��ՈPe��.�qeL 5&|���K�%0-�5Ցۺ��� z,; ��E(�N�EZ�7Ri��8 �����P�m�R�e4����Pao�
s��Z���%��&���>+�i�NH�vAb�+���Ec�!�8��c����~0-��a�?*YV���2}	�G�G�<(}QٱoIA)���(B���Y1��$������<�>]��\�.��p�O�}o
46,�N�G2`7�	��r�,��1�����R5�iT���%aS�,z�
>����,r�4t�a�:#NJ���WO m��x4DC�6�������s�C�J#�Ot!l�~�)�KU4d�o��e�ö�8�X'r*W�`��kJ�Oc�*��XN����3�͡,�
U�������6%F�+�|�����f��c�=w}�9�4���ns{KX�[��`m����9��ܙI�"G+�:]lxv
M�2&
 je@04�& �PM<	��XcB�	�΄�g���:F(sG[XR润0lEгp�9�,�Osʔi�aC��ۣ�;�mӈ�i*�J�4q�2e����0�5����e�cRlߦܿ���]�������y���I�4��Xo���9rrN�*�0���ll	�V�_KX�aS�I�����C�	���� ��L��=�������	�J��q��y,'غ����ؑ@�J��9惀��8J�&���Hg465��I�I���\|]�F��>��`$g&���u͵(g�W����"�F�󐖑������&�M�V^}O�3׆X��<�a���h{��:�,�&	0�wCP[��s���������Ǘ1�d#���'Q��*�.� �ϣ�x	̹_��W�K��a٘��}`ќ��TX���R%�);�2
�3���@�n�ʎ+㼽W*	��pe�����K����̹���.D�\)�d>��<�e!�%,���p5�[�M�^o��Q�n���g�H=���q|�~k��J%ׁB5_�	��1eЖ�������9�L;�� �l$[�\�F-�p���W}��~��͏��>��x���a�" j��k֕s���j%?A*���-H�jD�Xr��Q�ڎ6��o��&|�����T/��5�FBc3���0�o�4m�:�J�$ت�Մ�z@��p'uu����}
>{��K���>:����}h;ӇG(��r���~��l��쫂`X.z@�Mg{ƃ���,ʲ�߯��@ۅ~��� yٮ�DJ7�Q�CДmN�+�R5����]�n�P.z�0FP����[�6�i�K��e�w��aQ��J޸��6v�8���kj����z���g�X���x�����l��W��h{Ӧ_$dN�^� �����4�ypZ�/�S�O�6�u�ܫ;R/����(�3��;P���`�S�VD w�� |�_A��gS`M����H�_Y�d��b�ڡ,W??��/��엗p拋���v?9�"���u���-V<��-˳�)���xƻsLڭ��q§hD��n*����}ڱԈ��
@	��qGh��A���RSưNA�!����YA*��� TW�^z��^h��_�W>g�_"ӝ#��$8P>'{��gD��IL���@�yOt :tsR��
@'	���^��s?�� T����y��s8��y�x�����l��- ���$�Յ���T�T��d�Zy���'�8��E<��'��}���ۈ�����.'��Q��OD�@;�g&Q�܊��J��`px�Aq�E���A�LH�CjJ�*;PR܈��.<L�aQ)���D$A�HP4"�2ؙ����'�[�����p��-,��\�v������qL���_�����>��s47�#.6)��!4��bvj���"ܤf�c�Dja!�j�P�"!�|9��axfo�M�>���N$�c3ʑ�S������"��]�7����_�A����A�5��XI�30{7�g�a{�J�s��Ǚ�����5 *�#O�P�O��zj���N��&Xʽ_�P²�B���o���{��@�}H����
�ҠO&�@c{�	��J���X���(�Lb(�&@J��3>(����&$�Ѡ�2W jG#���Pc�&p�P �1T�s,F�x9r��Q@�@�����nؓD�C�2�Np�4d�JP���	|��#���_��	�\^Da]"�R=�w���(��;�A �$|:�F���ٜ�4�5eã5��
Ǻر������ jW��XTi!�"� ��c�oK��m8��"Cʄ2/�'��þ�N�p+��g�?|r}��h�iT�7"c�l�� {�.3�m��c�l_[d��#=��	~(�BAF 23�"%�(��G^t��G\r>�G���q��X��	���<���	��~0���Ԩ�8�JC|��ywd�����E�$����� TBpeP�~ڱ�
�ڏe�z�������9S������WI��_�єes�Ƹ��x/�F�K�~* m�x@�h���Dh$0Z)0��'�<?��w����8�������}g�gQuq�7�<�̍v�z�k"a�}YU�`���v	�pXW��z�ee�('no_c]����J8���p�!�YN��1���)a��Vf�%|��X�,�:3B���9�͡�d=c蹙d͠�I �&��P^\�d������(^H=g���S[�-�cee[+8�l��&3X�X�Fsnk�d#gs�p�����=W�y�<Y��cxJ��1���A-Y��0�`c	�Қ��1"M	���=�<� �>�3�VF0�Ѓ�� ������q4����l�alm sk�����5aݒ���V�hK뀬�,�=����ɘ���bB��X��r)���ʚ�u�����l,x�(��v��#a���^������xFܔ܏��㨇�^�8��� U'��Bdr0���?Y��p�K6��1���@vAS�p,��f���la����pX����2+��Y�g(��9~��3k�g�V���P�Բ/�G�J3�1^���"��/H1�o��@J��p�&ߕ�|~;3���ö=�����/ݹ����t%��t�I��D0D�s4�+��>ف�?��l��~P�R�*��^�!\� zd�G�K�'TBr�XL�<gJp���IY.ő�R�=2]F�,��0�;U	߱2���&��z</c �CӮ4�	5�N��@ �<� ��(��N-�2`֞��h^��[?x��z7?xcg��_� k��\��4*ƍ��%|:6���!u�3�Hy�m?7��7	7f�qe��9�`����B�@��g��!t^��x@��*8����˃J-��H 0�l>ׇ�ˣ�2�������E]���y�O�T ���(�Oٿ�m��0��o7�f��<�H�S��m<�������s}LyB%���
lV��:��t�����ܧ��~�o��艚�e���j|����&�I{��u�dE���|q�/$��>N|@���)�~HP�h_i�P��mD�th��)�O��pW>>��/�c�Әy��`G ����"���I)�I��2W�4z�x��/��:B[�]�=�`�'le*Ԕ�~[ƕn�F�� �=�l{__�����K���+�z�&.��:���6n��;���p���q��wh���[,o��n��.���&.~}翺��?����|�K8������f"�f�砼�<	7ֈ����iX�!����NB�0�Z��		~b�J*�/M|	�W	U�IB��y����:)O�� P�a�m�A�w ���O�ҧ�q��l?�,�����>����1� t�L�2�[tH �� &�c�@�z �!��s*��/@�@/�Ѕ�+�$p�� ����y@B��4�tU=@�2��	9��I��?�ݟ�E�B���p�Fd~�2��]S���x��Q\ӄ�a�m�CJz	�' H���D��XDGf 1.Q�i��r����8D�:	��"�$�����X9���w����1	��k��ǟ��<���z�F0N��fÞ�Ʃ3������|DG�#>.	�I�(/�CO�Z{��& Z���tD'����YR���4����������C���y���6$gU 9�	�e�OGhFZ��u��޸���I��ԩq�G
��[���^\��;8��M��Ψ��;��b�#³��}��Z �zoS�e���+����������5��m���� T��%�z0GX�egU��q�$��ā4$�F5�O�xvzi}��Ha�+ ��x�@��P�wc��೦�KB$ �������!ׄF�k�b	���EH-F�d9rg�Q�X���6§�e&�Xx?ϰ�0��1��	H"��O����+��?��7?�G\G�h%�g�-���Qp/��+�V�
	�M�KU�(���@	�.���(Ӵ$k@�jK�Ԫ:�	� 5��eJ젌%Q��2��Jy�>}ʠ�PZ@��!Xy�e��6o�x��ԇ`���z�5�n�v����O��,q4�AA��őxW�f�#�8�!�T���(\+����:��#��@�W�����g�Z�WᲞ���AU���������<���eajBu��-�p�L�s��em� �}?�sP��t��:������	��3rl����O�N��p���i �1�,�h4<��f�Oʨ9M�
>�l�ʺBh� �xEc�GԸ�pJ�Ӏ`h�Ҿ+As�h����onb�׏���������yt�w��`��qt(�m#zż�U c�	���3%�İ���UX��|.�i�/�ݠjCx3"��9�0���LL�aan���0�4���˂@fM��|	d�V�XG9�0�	zЋt�A�3���`���$o�'��"�f1^0�~60r����1-�`d�s��� ��
��������0�&�,�Y��0�����Y�/,ӎ�<�p�����6���n�s� T
0rV&ܷ�)=#ʜ���x���� ��}��C��l��3���i&C�?,�x�g���!�Z��,2�������F077V�Yie�w��򾒩�~�τY�L�����ׂ�7�~Y���>�31�5�����y^ry~���k#�<��'� �k�7��
�G����hx��[�qX�y����>��^�0����;���fnV���Qg�#w��~���y$,��Q��g���F���9�7��<SF%2ƛ���(Ób���l�g�O�R�6U[�?���#@:J݆����7�����?q$,r}�zs��Cx���s���F�weFup��@�N+b���T	Ϲ�K�-!T��^��QIPT��|xO�KƁB�W��X�#3�8�P���g4�p�� Bh�bfa+���g�gT��h!��E
��g��6YK��FmI0�;ǔ}� �y,��P3���M�!)u jB�4bk&PI�u�;�n��v�)���C�����&�+y؟Xp-V���[6�O�&���ʑ�І�Y�X5�fP�ځ擃�D���/� 5�)^�Za��^��
B��:ro�oL���Z/(鹿h��At^#�RC7dz	�,��.�?>գ �Q2���P¢�_���
�Vl7��[�fh�~r+�)��z��{�����\�)�K^B�<+p�d��$N��2�i��%���q��n��W�% ������ ���3�fɃ"94��"AFBpw	W'?>�S���g����a�S2�g��J()Ӯh�}��Џ�����8M����>�Մ㾷N�Y�����
@%$T>�� "��^	��=�`�� �u��=oO��m�;��#���7N��~ok<�s?��7�6n��>���^C��~T�6���:������EVw�j�\����T�tf���i�x�gjѼҊΝ��b��������Y\��
.�����X�}�����I���<$5�6A�H���u *^R�XP���%[���A��x��- ;@Ŀi!�u ��, :���V�@o� �.~r'���&���h�~�_� (���7�1F�|��1� t�� Ưa����T%��U����������=��2��%d�1���t��$�V S��FJ�Խ
�]S *����o�tV�nc���?8��?z7�S����ɎBDn<bRQ�\��Q� a�����?���:�E����a�I�'!X����#"�����
�#x�� !6�q
���_�Sz��l�����^�F%!(4�'��~�����72���^�N����¥k��mDNN*+j�������g�c�w
���HK�GVV	�1���t$dd#����m�����X�;�҆vd�!��I�HϭEZ~�K��2:�7o��[�<����N�T �5��y9����.���>Ǚ/�k�� �nK�74��>\-�N�%8-J� T�S�~��O(�Rƀn|�{F���
@_A�4!��R*֫	u���L$�BӑĎ2��};<��\��B��m6�{2�R�%Z2U��*�.0�)�1�tI������� jaN���H�W�?��_����ՠh�U[2���=�G��q��F��!vz��hJ@LS����5߁�wN��?|������+h�-��<2}�U	��H���a�\7	�%|�:���5!�\�w-�:T>�bT(�5K��(�0���^Z~�d,��R%�R�)e\��I�1���}aP�S�Q�?��`T��b/8��>�v)NpHr�S�\S\�����ABz�'��CM0��	�<��fUGÒ2�%4�N�@��z�� �V��`ϛ�bT���]��@�������B_�fe�0�$DE��ܐ���<x��tlK�c;%p	�=��P���p��O�1��4R)��l5EC���M���=��5��PD�4 x���,�iS"�2�
@5 *��- �k��>԰��ښ��Ԅ�8��x�	LV����o���^�Ʒa�x���e�,U��T������ʵ��-��|�".���Ib*���?%tub���4��}��a�� X�����{(PbOh�#l
�9����aF�y;�$�W�9��[�ZY�*�aS
;��M1pi��k�\	�N�{՚7^?���L&ds^r ȝ���1Ý`�����e��#S3^���>s���.��t<g�ep�0ɕ.�����U��3���b�}��(/�gU�,��ҘB�/��{(�#2wl
\F2�X��
٬F�N=��+�G�ߙ�ͦ0�	I�x���#��=�Ֆ�ǆX��EV\&�YJ���oa�-PF�1�y&�dla#k}X�w�P���+w�F�y�afB�q�!�(�raN`7&�����,= V��`���P���2;�9A�)`]q�Zg�����H��}��~�#��<a� �B���T��>�z|��e�������V��U��p�B`(�r�J��uq ��.㾌J�ި��Yߋ�I�l�OW�W�{\�X)�������`�"pڗ;��mɰ�w-�>0���^M((��,���!� ,�P��$�\*S��%#��Aq� �|/���w��,�A�>r���U�zl�us��_m�љ
�2o�7ԋ �5L��͇Sw.|h|�9���>��AO���;Ôω��P��<����w&��#	�P��$D�d�ԓK����o��_� C�S�໫$�|-r	�f�)�m仲9Ǉ*�F ͜kA*4��+���U�@ͧ���`���6��W�����$

hܞ��;K�,�u}TAh��!�zcZ��+ ����%�W�BOv��u�W��
��*	��P�ƺ�v^�"��s�-��~G�j�+��O�]@UBo+�s*a�g�*o�k ��\�ӆ)��d���������g2}
m�'����e:�����O�F���~vAA��bW�K�խ�ģJ����n`N�qF�<�r� ;������m<�/�|��D��R�<�fK�T`J �~{=�>h?T���2�˅�����y���6�*6�D�����y���}�3��man�P[X���m5oC����� �|׋�Xg�k���p��k�3\���`�wY�۶Z1ss�ˬ ��N���k,���{�*���d��=B�2Ż��mu�J���e��� ���M��I��߂P�7��ȵ��@lRr��nj���� J�$8�@/||�,wo�|-�v����Q�ht�1��I��] ze ��0�:�'>���.�S T���̫1�_�%\\���ب��D�7q������}켷��������-��p;�PK�%���x5Yq��i�����|N( ���럜P��B��HJ����j��2^p��p[*^Ѓ������/J�%���'��x~Ovp�S>t��!o�Ή����GD~<�KҐZ����6t��P���Jĥ����X;��d�%(�	�G0v<��
<�>>6!���B@P�G�q��C�y�U���?#3����ԅ��*(B{o?>��s������'(+�FMM�ں��NpJJGTx
Ξ���o�8��� ܤxS�'���
�uM(�w�&����G8w�6��\�Č
ĥ�"3�ye�(�����&.����:�fzQ:J��+ETc"�����]ƃ�x�;�g�������O��ʋ5�7?�S���1���RP�T��� p>O5��@�@� ������pKy;<�8Pm;����}��'�f�и�$���"��N��v�i9 ��D_4�\%qY/ZDHL ��z���JVL�N^�S`i� �LꭌaI �d�$�/���K ��?��d�!�l�T9��Q�܀�v4��G���zL�'{Q�T���`ǝؔ���6��~��#��wq��6
���×f�����Q��0�>])~v.���@gu2+i�S���p��j�a_{§@�ue�PK��cmV!����qP�e4�"�e�z�rQ Lh@���hV�ð:��a���a���Dk\���#�ࣰ�dY�dOP��%�ԇ¬�8L��`Z˲.� FX$T�.��� �G�������DT����( �Ȱ�F�!Tr�"1`��?�[h<�$�Iy(�%	e����lK�ow6��25P�� �:��aX��t"x:M��e� �E���\B�L�bT� Ԡ&��3��)
F���$��4Ra��j��Q�9��O%� �^K��b S�3�AmH��TNJ� j^��/���# 
T���pΎX��07�AnH�O�Q�LS@c]��eJ/��Ђ��e�|�P�J�,��	�/�X��m��"\4����0�F��0M�E�����m�Z���]hۄq=���%���k���14~�`�ǞD��~8���L�p��^���ö{��9� `���~,�c��LXNry:V��$��,�fC���r� NK%p�.�AҼ!
z��I�u����6�!y�m`� C�pZ*��b1��a9���t��f�L4���,��ȼ�l;�Ype:�C���k��k�kB���c�#:Y�-	����$�zʋp����(����A��������|��J�t�%����y��~,�xa0J��]Q�����K{�O;�K��8رmڱMڲ�۱MZ5Fì6��1L��P	�3g^ʌϜEE�M�|OD���.�X϶j.��w�$����2��Q�����T�w!T��Ϯ h5�)˔!���5����$�vݩ�����Ʉ�a� �1R��b�i�s�J�s%�9¾��0G 5�3f��k*�b!�Js�~�3�{�uy1�ck5�^ ��q�%*+�4`���U�y����#�[(�qB豹R�O��t����2�g9|�<	�E�]�_(�Q��Uyi���u2M�EW:Lړa�A(d�hޛ�%�b ���e�)�ٟ+��5����	0nK�5��ޑ��q���)�������+�_^���e����k�khٞ��4���'5�!l�
i�Ȓq�Т�fT�u�iw ]��yaTy65��!���ө>k��*�[/���B�x?��&ݙE��)��9����W��M����Ͼ+��i�^���)L�A}o�:��i �������[*cMu�)�+@*c@$6U���}j�$ϧ҅>�]WG��T�U�>%ėҍ��E�����T+�L;F�N��.a��sX�hK�����=�=F�Y�pE2C�Lò��6���΋}���s8���?���$%���D-\�(����3GM=^�����ƁҖ�#؈T�G`S֋u�*�$ *��~+0*�������z�NL	8��5B�����K?�I.���7f�5V�`>������*���.����G�;|�=냣�o��"�p<��Ѿ���u�����Jޑp!�;�� �j� s�G�@Z�|>g}���߼��9\��M�|~F���k �G��!	��$L
T�<��%ੲ�R��W�d�M"B%���	�����T�e\�Pٖ|�
B5 *0�AqY�_�;���'�ܛ�؝IL�|��\H��/����38��,V�j t��:��ѱ϶J ����m��	ޓqLݚ�8A}��"����J��#��b����CX �#��}���s�kB'%P��c@@e��36�w��J8������y��<��V	����.�)S���o�)(��/�	^������d��lW���)�k����W^P�PIBC��t�=J��f(�V�9%�>�pk�k[�C��dG�9����H��E!�8�EIȮ/B�p7Z���>4���aW5!-��q9��LGD�&�6<,�\�1�)���$^B�p<,�~8���N�4v +��	��;�#�(�����y������o������#����agw_�K�p�޻��mDXh4�D�0�}ӈ�HEqQ-j�ڑ�&��	����u�Ե���'N]���
��#|&fV!9�
I\�,j@b^%R�k�8×��(jf:�;P���d��Ū�Ww��]<��g���7q�����)lzB~K �{��{AP|.��T����m����9E0�y*���=��b_yB��a�V ������d��҇�]�2;���dDw%�1��~{ �J$l&:�����NV�S 4M<��RT�,ʣ���@���z�N#�ᔩVL�t"�@-�d��@-��(sc�j=�	���)G_�94
kP�J �nc�֫�*cNX֞�@�D	B�а�h4�����������۸{k��YJ�W��i�{�«(~��N�we<��Z��x8W$��u.5,���D9�\�4bm	���̸"K��E%A���a�р3��xX&�Uc%xr�U"�}�B5�	aS���#��pj�S�ڣJƔa�Bˆ@�L,J�uzuߕ�E�\6���$|>E\6Љ cXM��D�QQ�J����'���Ӵ2��7������ڜ��4@%׽-��P��Tm.u��4���l5�3|�n�=�vՑ0�0�:�XHv[J2݊$鐡��>%�V�z/E�m���)��xCu2!��L�u�mRֆ+cܨ&�`�5�yO�@)	��>�Ӏ����$q���WJ�!E�݊GJ<S������,��aUkʆ cS��p�ϧ�0Y��Q�}��)���ү�~#ۀNMT3�ζ��.Bvw8�{"a���T����}1������=�
��d�$È2M��X2�D�4AMRS���:j���\6l��Z��[u8B�m2(��jX���p2�SЛ�)����u���)�Ӑ2{%��$B1��mȅ�+��>�p'0��	�Cy&|�	O�v���%��1�>�Y*y�с|U(R
����[ 7����p���G]2��S����wK2<��$�����Ƕ�6o�w�Y7ϻ+z�1���P��0���vá��{#ϳ<��|��\�U�����ԫ����V�f2L@��Q9��C��0z� ��@�]��Z�Wm�#aٙ�lxO��]�E�f3���v·�P����c_�3��9p*Trd�!ˌ���D��¨)�MQ��l�4-�	M?ۏ�k�*$7h�~Kj*&ϥr������XO§�h�����\ߩB�Q�SE |*M�(，��/��d�����.�+�Y�C���y��
@;	��#-�?Z�oT JP��U�)c=�H�^Q��Ÿ+�sɲ�϶Ӻ7���?�G?ŗ��7v���wJ�5_��ܦ!��I��M�O{�Gk�6��>��c5(�%p�v��� ��it_^{P�<,�#܉�����G�W4��,�" i?�}g����u��A@%��'T��7���������}��KlT�݈B��q����RN��SJ�)�)�)�١����W�*c<��)YoeYBu%#��3*r+v	���T�.ta���9m0j�����)���?���P�~Ҟ ��+N���{أ�O ����)PP���\���Ƣd�}��4��O�tI�z�8BuI�t�	��$Ñ1�:鼡R/ +Ӝ��`۟���k8M��m��5Ѱ�w�E�5,�[Ӧ��C���'��3L�"����-\d^j/+8yX��������aeo'Sغ���3��y�>���0/��xR �(�8/�G9�,���z����W��1��s�O�ƃ�z��~�
Y�;����U]IF4(�\oM���8�6d�����g����*�8 �0��) *ЩIH�P�f��:�<(�=����HR�{<W���{`�E���;*���+ ���\�Cש��@��Q��Y��=�	>Oc�2t���򀮾�����a�Л��b� :qmX����i<�ߜ�H�Z�7�4���חp��K/ǀJ�γ=���V� �!��<\��:��%W �u ���Ë��|'>���';��t��d;�f��J����#��&k��i;D���M,�!Y{��s�\�ÿ~�\��wJ �R�"�0S���B���`luM�������MTnUH.�cA�8���d�V#7�I)2K�%,6�i9�.(CBj6��D+�
GAi5j�:�ٯ�Y�Ԃ�|���?�'���Bw� z���٧_��?�fg�iNDvfF�Q\X���,�T!3��Ж�^�w�������Y���>ڇ�Q�6�����n#&%Qi�������
���Q7ߍ�zD7�"�-]g���/���/n��O���O����+�\�`˼OK�O�2W+%:��|N<���{�#M��:��H��@�@��P�� t�`*���� �Jn�H&4��I����Z U�D;�dh2;�v��P)5�5�Z8Q�ԶLX�[A� jB ��%2�����������ʂklg
�?�7d ���T)
�P�"�?e��v4�x��N5��n��"j<�5�0r�4���2>��.>{��'�v�� ����9�.Y��Y��xF���)*��\�(�Ѫ��$*9U���r %tڔG��P�� j�:�Jr+Up�3�1i�R��J��!e���$lV�g�h�<��S*c8œ��x�h�l�jdH�hJ��^��-=�?@Cx�ie!�i���)�~�$Db�;w��S�	וF�ˀxRRaן�ƀ�$D:�A�Bf�`A#UBbMk��B���$p���4��C: %p�'S+=Q!��ڹeHq�A��� ��(�v�-��Fnh0ׇ����஌z�'T�I��UJ_W/�y@��o�´:f�EU۝Ffe�qx����,T[ѯe�4l�l�}�J���] ��%T��m� j�A�o�&��E@(��<��t�,��d"zC��^�^�^W��eH P�cI�Sj��y��O@ԟ$��Ӹ_ʅ�d:�S�0����T)Y�<(��>Ʃ1��3�pj�S@T�To��ͥ�p%fE��,��j!�V�`�Q
��2س�_-�A�e�nT�Zv]/��J	���/��q�6s��ʁ�T.�
a;�;�a:����$�|}�Ҿ��޵�M�E�O����K�QG�O(�����R�ϥN��T *�|>,����{Ő0g$�)�>)P��U�x@e�>UI ��(=B�TڸqG,�S	\Y|6	�>���<8��p`����z��3A�Y�o��Ep$ �y��}9��{��5 jD �h�Q�+mڝ�M9Ճ�S�]o��L1\&��1W�#�5�#|�Ovٿ���i8���σ7AT%&"��N�^�/"�k��'�qt��e%<�!�����-��SAh7�hGL�4^P��t5.TA(%Q��5vӒ}��Ԭ/F=)0��ͤG�l��� �ӕ���<�����_���콱��^�\��� ��'�P�X���D��>�P0ӊ"�h�\3��:�yv#o,����w����$j"��I�m��1��1�Bq�2��� ���0�E���)cB�*���7I��ܯxV.d�h�xA	�:ϧJP$c<	���T��j��R'0*�iZtc@����u��I� m�1��Z���E�
=٤�N�������OOb�jY�Sʕ$*m��	�O%�v��u�tW%!�%x�#F T�T�������6>:��w��\rqlb���u
X
`
\�<m:�<��,Pt0TT<t��.�4Ɋ�	-kOO@O�8��3(�����`x$z�>����PG�;����^6�q���lB����V,�l��n�#�<�����#8�/?g��oz�7���`jkK����
�>�p?��`W�n�c=��
7�b,��!f�JsC����"]�9h��6f�Ӧ�G�&`�xQ	uO�$:���������e��,���+o�,k��A��ɷ$����D���?�	����a�>����<�q��%��Wy/Ρ��(�7:�sv�7���ޜRYpe�ɛ������g�*��(A\Bp%��#*�
�=�����I�TP.+�T:�������s	翺��N) �x~�	�j�
@�$o`�!��M���P)y!^������}��@���:M�&��
��f1�d���|W�v��&�8d��7��~�o�[�6&.��hn\�\�2�/���x�6�w~�5�����x���;����G�,Bt�4<�)H�.Gf^��%��mݨ�o&h�#��!�qJ�Y���e��[����6�P�Є��	ܺ��N����
��~b}��h�
�Q���
4��!?�����|Ԡ �����*�L�R���!,��ca�,�G���,F'�\P����m-b��	�m��|���y��C�v�}���s��t;_�|���s��
xmx�@��S��5c?�xD*����cA�%¨�oi2� ��䪐[§Z&���,���x�`O�^<�I�z�����9j9�OS����|W.l�o�3kB���P��@M	�&
@���7o��˵(_gg�%�Mw����Vo��vv�R�<�G �±�P�������O����pq
�������5�Ni�p�<
�?�g�+aԵ8n�1�츄ѪD�V��MBp+b���8�>u ��Ԍ@yX���<(�x* =���҈0��J)�x%峉VjM�z+�4���r{HT�3d�:1n�R�*�R]�� ���k��k�G8��9� Ԫ.vM	�!��WIxraY�>�4�@��ԑ��ou �:�AÕ z(��h<i@_���`y��*BaA�� (ᐥ�fE��P-��1�N�FA�/j'��P:�+}��e���D�i#hv��o'<4Қ�����j�=^c�+��I<�/��S` �%�+��]	�^�1p�ph�'��-`�>>��V�<u�k���A ��>�"a<�d8��=�~����EJ	�I�!¾,�F��	0!�SF
H	��F�C�	��D��ىd�S�0�J��4%%��B�`h��A O��꼣S�L2��y���<K���Le?�<�%@+��s0�&<��y.�"�^U��e_���k��}��k�ڐ��H����z�����u�ݴE����
t��k��J: %���F��	ea0n
%�	����6%�?�$�^B���C��>���2��{Bڤ��H#BH��xS|W�T_ P<�u��M0j��I7�+%0j���@�2;�a�@��	�E/Co��#*С��ekB[�l��^#�N�a�-��GP-���cpc˾ y��'�pt���ڬǑU£L�4S �bx��'r	����jA�gL$�I��k�S�82U�ƀ:��\��r8����� mM�i{
�;%K��&�}��R����#��l�~U��C�~L؏���¯'�k���O>�/��x��C�{v�����4N/���4J��1~�$JVq�19�-(��@�R/jWzаNH�@�%�B.������:�/���
J� ���P���/c�u�?;�Bo6'�ZTu�7���_G�e�܏ ����O@Te�%�ʲ�I��˩�M�z����Z5��9@�\<����� j�g�U��#�ی��Ԝ�My���F1��
V>"8~�����$��H�mH��U�ҫ��W�n�9A���'�C�^$6���
�S4���6%��4%���#�.��M[|���y	���0x�΃�$�[/c@�n��I���2�n."�����L���.p	��s���`�f3#�����6�GGs�;Y(Y������q��*Bm]9��+P����,�\*�(�I�p�r�$�3҃�	��TF�z�$���|B]q4�Ǔ����PkX1�]�9��O��5������_�W�s�'���Pc����)��P^W�E)85��%�,!�: ���w@�:xO^�J�o��	�N>��~Fy@'����q�˛�z^e�U z��9?���Ԭ��i��|@�o�(� ���Әd��;d�G�{k�7ض�) �~cL��>#���O§�=A ��J@���3_By�}yQ5Nɀ+a�{�ƙ	���������&��c��M�>^�	����B(�F�] �\�P>4;����g�
6�>�Vਜ਼~��� "�#���LM�&/>���?�����O��_>���<���5�4'�+���G]���T������Z���"�D���X��&�������u�d�����x$f#� XZU�����{��N�L��ENa)�{��Շ��z��c��)�W\���v�,,�$�N����4:�{0�?��df�B� QI�y�H+ArB�	��%(̭��QUو�V�$�:1���͋�1�����a�t����=��A�j
Gj��]���T.6a��)���w�֟���?��S?:�_�a�],��,�:/<]¢L��r��\�\���`L'�V��O�nl�@��'	�/�x�Ք+�t�*sʘP)%T{��h)R���!I<�z ��X48@��⺹;��!¨�.�ɭ���o�S�9T��4���\+K�kbo�X?ī�2��k����[ͨە����0�~��2��� �x���,G�`��=�gO��Ǘ��V�#�4)I8Z���
B��ny��(
�$%�\J������,1p�I�CY�Q��$�UD+ =�V�P���O��	�5��'ۛ��(PI<��&�n�yu0�k	�4*���)��?��)	�5����.)#�.e@�s�?��xXD��N�O��emli�6�*�q)��;��X���#�F���G{�<�Z�iXRi�RC�t�Q;��Iv���#�"Vܿe=�_J�4�B���S��,�y@	�"�O�T���)�'T��Br��k%8��)����@�x/�h�
8@Ux�k$�z���k)�kuR`��1�\ �(�42������W^1��&x
�����l�~
̴��@+�VBE��v���#�O��#pJiD�4�W2�"��Qü�ü���.J�� �J�����'��h:����N����ws<It:�)��D%C�@��S�kd@@�Ȥ�oc�d��a)���ހ *^SFG}�V���!�\�����r}FxFy^eyP�<��1�f�w^c^;�>Be�K��f;c�`�i�5?$�>����I ��6� �0�H�J�o�߼����k��Y_�}�t��= �*�����(ɀ�xNu�lC��H@M�x_)�N���X��g:s�8���,��u�χ}_��raݓ��,\:�:R̽@�8��P�&^k��ξ)e�Uw�{u�[M8�Z�#kU ���6#�L�7� ���y*�g2�P��b���$ *TӰ�����BAh�d�����o/�@�uW�
/���xAB%WƅZ�Q�Gm��H�����~S :��}��(�Gۉ!���g�◟�ѳ����'���������3���'���c<��b��&��J�7҄�4Hi��n�v��uN2���$�?�J���+�*�V�{�X
8��h�N���}���%�v	��M�� Z�˘P	�Ս�2�<�2�S<��O��.26T�V�SJ	� �����@%�V<��]W��_�L�"�<e�`�xAB��*��Ps�0p�}o�+�\���,m[���������;ئ]}ⳓ��x�`�� t�C��3������t�%�ξ�����_����J[
@�*!�j+��:��e �gLd�g]�|���+��O����I���!�v�g�'<b����#����=�l+{C���^�ӎ�io;����JRg�uA��QP����df���eiyj�+��ٌ��5\�~��1>?���^tu#%-n.�������m[W38x�Í��o�#�b=p<�~	�8�推�`�����gq��q���y�OҦ]Ն�ʵ�� J�9>��
l��T�����
�_J��;�a}gco�`�`<IH�~kVy@e�x@7����}��XSI�:O�~�v�.5�����C;����j� �̽%,=������o�c� *!�s�&� Yp���<	�޸��4N6��OaO�~%!���4,�eP6Pɂ���N��* %|�$��t���ɖʂ{���������������{��|r�|8v>'x~�	��%����N<��* �$�L|枮�8'�pm��O�����?�������3W��恀,_�W� �F{lI<2jr�8ҁ��1t�Ϣ���yH/�C�8����ΡYT4� .��)y�.�A~i%��=���oiGAiS&�.Eg� �K���i�7�;���,���bX��v`p�=�� ��K�<��	MK.B*�����2d��,�Ey���mEyC�:�����Ao�pw�/��'1�=�ѓS��F�l��Ӛ��uOO��_�����˿��?����v���	���%�N^�y^���y��Y�_��C��)�9��4�5�5�M@$ :�˒�z�K��K/�y��x��S�vUQ���E�Fn��x��C�H�a�D ���G�(q��E�	�DPv�IM)�;����sM�A�P��yG��X�6���L)�c+��Ŕ�De��T3�� ���6֖0�0���9�� �9Y����[�6�r�	�'��(����=�܆�����#�@|��Ր����|x\��ϯ�ݷN��+�|a�VF#��,�`���� ��)/�Kע��FÉ@jKHu�(�ա�PZ��F�QE�w��V��HBn�)A�0�J�Y�K��KÌۚZ��f%.k<� 5�hM���Ti<���0���k�%I���% �Bu_�R�z~�6�ۈ�I���Q�Gg��qj �0[���q�+ ����kQ���X�KS"�����Uc��i���B{��O�U�  ��IDATgߛBc�:Hcm$S���x4�/����ݶ%	�[c�O��OO� T��Z 5l#ȴ'à�����գ��zP���~>".��`��[���7§�^5	��8;M��:��LS��+�ԉ�����s�NPJ_�ke�6 ����4��m���S��z��<Ƕ���������+B�@�
i/� c?��B��'"|���W��xL-�*��$�<�e,�K�� �
��y.�y��[)�<*�F��c�x<������\n@��� ,����#28�>�y�fTs�9�oF�5M"8��~�p�ϖ%	%f��	�F��%��p&<?��9?��2�݄��P���ϖ��`;��튀~7!_ ��`wD�π>W��: ���G��K�t�c��m����>��-5����Kvk�3J�����Y�2t���k5�i@�4l��a#ϕ�%¡Q���׆}���!6�C�{�`��Ϫ�x1�G
�<�ö/��a՟CX� ����y4�Jc�k��]��� ��L@o&�R�������i�㳯��W_��~���7�^��rm�"�R?rh�Ŝj��l<��O/¨$'�*D�l)f��?MM��o�n|y�/;6[����i	l����:W��/cX%1P*!4��ʮt�4������z��̅�H��P�
��u�;-�L*N���_��ß��/��S|��C���M�{����.�������!n~� kw.�j������F�lm�v4���e��4|�Ώ�?�$!:(�����]$�^D��.t�E��!T쵠B���AUI���V�{�^�񼭲ޖ�ԡ����"$ܘ"���f�������I��DG26T<�
D	���2��� ,������U���qeL)Sy;��A�� �̸�Y(�#��9W�nA��64]����	,}���˳���h�f%�ЋMl:O��ߜ��秱��	5���GЏ@	��ݏ�N�)|�C�\���,2�	���i�풄h� *	��d����M?B���;�1 ���u��}�,�n����>G�\��]��3�&�q,-ޱ�pw������ưt0"|�����F��1����F��p��t9�����1aHKK@`�?BB�"+'}�]X�Z���2�sLizu�g�p��Y�^����:��QQS���p�x:��ڀ�����a�d {wS8�Z  �QyA<oo��:"�*�s��g\!�B��2��0|��d��w �v>�iH�)����M�ɵ&���k2���;�aX<�ߖ$'�ioJ�V�u�=�+tH��ޥnO���dW��`��SX#�ν���Sl�{�h��A�~��b���n�)Ȕ$D��Eƺ��e��<֛�6���X|kK�\�]�ίNaK<�_&�<�S�\����W���y�>O~~V5�u^��wW��h���a��I�?a����h;�U�-6�R�:/�:/�x@y�t��:�JPċ��|{�`�*�7XJȥx�4�)q�">H��P�r+�e��e��g�yg��~�˼R��"Y��V�'p���	��?���c��V�H�q"�4q�I��MDZ[6��G�}�V/^AVM+��S���,�	��3(mnGjQ�YV5��������r�t�qWW���]��fC�/�Bn^A�CS�*S��N�ba� N(�^XRS��t��g`M�݈�MCbB�SK��X���r��)%�%��g#/�Y��Ȫ*B�p'6o�㽸��'1}�$zN/��/���MW ��EK-��������g���wp�ױ����bKo`��ꮣ���G4�� *�=�|8�I��i�*-(��{O�v����1n?N���1&�.bL�\��(\)C�p�	�q����KA��~Q:�5R�O�`��|N`�P��ڙ����%x���L3��L5`��w���
6���R�>��aik
s#X[�eI���n�G��U��ځ��*-W�t��A�jD�v3�����B;��KC��C�<���#��@�h�~�*�=����������*D|�1DU�!�.A�p�	�k�Q��t�9ׂ��8��!��
��^��E�J]�b�Lpu(��mY$�)��X��ü,�"&-]2.�J��UpY$=Y��B�����^3U�LߢƇ
�V
��'�@YŒ:�YdD��`�^!�j�!����D�<(�� `@��ք¤.��Jc��PY���i�ʲʐ)����������62�J>�oS|z���OC�'��)�,%{�n��Gr� YUGsa/c�d�V9��d�O��xX4�h���1:�bE�g]L[	O�l$�O��VBFcQg
��R! *!��=�E �d!&���@�B��#����8M�M��R}��T�����5:x���q��^]�^;�$ۨ&,��t��L�P�t����G����oK[�M6$�U�������� �n	9�%>�H I���IBk�5 �Bk�΃ ��q~_���II4 (��	{�A�[��/�{0�m�)8�K� *0{P��V'��w�ߪƺ��O)aU��j@�ry�ׯ�mF�������ƀP���+�K����F�J�	��&��&>��S���z];UmUڱd�%x4��0�v��C2�,��G,هX�XH��(_=�cK�aI�C͆�LM2�>w��3�/a��gO�(�S�I�δ�RB�ky^e��!��.7 n�1��*����JDl5��ZB$,W�l�.��X�Jh�<�7~��+��w��'���t1��qt�~\>2[���J�N�gB`�R�.�j�mG*l(�N�6�Ӟ@mO8��yMs��T��zb܎�9\.@�\B&��ז�j\��:�����=��ۏ����7p��{���?�
O�^C�� Jz�P5ֈ���L�;�D�m��G�Qt�F������"����\?Z�mW��|e��Pw���j�w��t�K��5��dJ()�	q���(ީG-���� �h�N����3=��iA3���8��$����[�g�&|W T�MWƙ�:�P�Q	���9*O����D/��
`juYoB���O	��e��r�)���f�_lGå��ì�����ck�[X�[.�J�퉏O�y,�/��G�j�O�VD���z�.>#`>]��{��c�u�hc?�X���E��=�=�h�d��F4A��m�������e#\M�{�-V�M�#(�\@��q�/�"�*�^�􃻟�	�V�V��� �Y��$�Z��6L���-nk;gB��-�\���u�\NKM@~^�Î���~�(,IEW=Ff{0�>���1L�L`��<6�n���hlEco#z'��3ދ��,X�������V�Z���m�l�삣	�8�rG}�����/�a��6���8!\���|I��R�\�C�\�h����m�m�e~G�gW	�kdK{X�)�>i���^����Fx_Gq���<�Oa����Lǰ�xK�@�z�v��<���a�����Aǉ4���y�B/t���oI2�)L.gޚ�ܽE�<��3�g1yc�oLa��fߘ��ݥ����ONc��M��[P��|�%��=&<J���i�PIB���l�����>�j����:���n.Ѓ�� t\`��2�D��De>Q��/N��oࣿ��37�ŗr`I0|s��xI���ߐ���
L���¹��CDV)�'�!��ie���+Ffy5�G�6<���)���wx�`9���u�4s��QU[���|�䠰� 9��(��S���ك��a��ۘ��Ne���~��zF��[���,�gҒK�*�T�,hN�3�� Z���L�g'�����{���L\�D��0��e�jn���T��c��K���/����	n��Ǹ��[
>7�~V>���X�D�u{�� *Z�p�g�j�r'@��~ �Hc����4�h�z��TM�1��@������)N�#�6ޱ��������d�u����L��b2���1,,	�F����0�3�G�?Rڊ�97B�Q�R���:Tnj��_z�|�鴳�:��7��FP�Mu�m�rZ3������7�޻l��P���[��� -���Dq���x��1�(\��N u/U�(WS��<�+$1Q,�ʢaWJ�,���[Pfl�f��� �H�S�>%Y�9�: =�%5��MJJ��R!��Q��E��A կ	���k �daU�AB͊�aV��t,P ��6�ޗGP�N��!1s5 :���x� �1Z2݊aߪ9�mF�>%9�I��0*5B�d�O���+jy���ݚI�E&��Pc>�Y��	4���WT`��@�T ���z�P�JX�N��Jbܿ�_Z���*֋'Y��X���P�j	��GT��f�-�ܪq�ܞ��	��2	�©�Sr��3��+B����I�T�NP-|��Pp�!p��� �aO��7�R���^��P	��~��P�OH��{�NB�@������k������o�9D�������a�A���;_I>u%0�`M��'��u ��dَϲ�P&���|�	����8I�N�-I����uh��
���96m�5��T���_�&��[��iF�r��T<�|g,��k��%�ʔN��|�>ݹ��h\���_(G���M�c$���Պ��5���p\��9Z�B��xn|�Hi�w���K�˼���pⱇ��1^��R�p_�U��E�Z��1���O��q��\y��=���_?���|�'?�����.��WQ8X���ZTL5�b�u+�7��B �>=��S�
>u *�6]B#���� .ʸ�Bߍ1�.:8�N��e�����L!�e�M������-��V;��~�������LH�����F���T@�Lt
��:�z�7T�AȔ�pY�'* �P~���yDu ��h9���[	ۢ6��S����T���32��W���!���*���*�o�T�[�.<!�>�>�[Q0�[~	����+
8B�h��t :Jf�+^6�} ����e,=�}���n̠t�Ǌ�`�ˣ6��������L3[s�VN��ӆP)���4�#
|�z;�����p�tV�O� /TV���a!G��j[K}x�����>~ΈO	�]����|�6a|uK{���^�!5?��h����+��m	�_;§���ehg3S8���7���A��ADQ(�*#��g���0��ۢ��~@�x���3�f��3,�B��O��>X%���΃z=���2�j�ۄ�㽛�~��@T t��)ާI��7F��dW�|g?�����b��.�@/΢k���V'ZNt��� F��c��B�{:E���3�J��k㘺>��s����.~ =��%�b��t���e	�}����O@w	���M� �H�+��E��N^�+��� =,�|��&�"*�t�$ $!��N������҇�X�hK�з~u7v�����)��T�8�M�T/)BTM,��Q�S���at�͢�w9u���!dU�#0>	Q�9���C��<z�f�7���C���id#421q	���Ejz:��PV]��Ih��f[O&f籶����]�������YW׎ؘt��d!#�� Z�tBhfr�S��+ �����t��$���
�7�p�ˇ>����^M5"��s"��V��N}yO�����o��3��������������b�pi<���>��} ��5�~���OwUۘ�=W��(5�{ 4�FA,��=���JQ�<(I4��
�~@�MW*��17o�a�
�����'�<׉�*�F��=�Tx���F_eS� �Z[���X�S�� d@�'P�\��U�~�+���Z�ۦГh;ߏ~>�|�3��a���lԎV��3x��:���S'PI!�.
���8Z������#�=^HP�� ��­ �0
��x���K�U�ñ4
�%��,K�a.�IX5-&|�,��BaUN��XZ
��ô�ZoUA(}���XT���t��a%�[ �`�!�$���� �ƵJ.�9eZ����#�>���?�Ϟ,x��i0��<)Ǒ8�~�<(�3��18W=��x@-��`ޔ��x�4A��e�Vx�^�� (۪	Ԅ�֨;���>u j$�)ڟcӲ�QCQ���-i�@z߂P�b�k���2�Ż��
qV����묫��}�1|	P@�ҫ�z6_�znO�4h��f�Ձ��Ӡ��SB?	�ݑ� BF�C����B
<��З�C T�	����h�K/A_+���j�/ O� ������~�wt㖿�W���t���>۵�u�N>O�>��u@�#�v'��/f�W�F�^�f,G�&���z}�@��UϞ<��|κ��DM��Ps�9K3��gٜ2�g�6
�}�H��FʙnD��Z�D �Ic�
��%��\��M�y"We��y@����;[��K�aVj�w�@h �1t�� Z��R���s̇�vY�׺� ����Ʀ=��Z��b8veæ-��pʇ�d)��
�9��Lx7%��D>�����+|��p����F�|j�ǭ��r��}k%ҩ��B��� w��(�b��L��$�����Z�5�Ϧ3?g�E���Q���z���0���h�;u(fy<�N5+�>ׁ*�b�U���]��!��l"������CC��Y�NBc,PeY��2�T@R�S7�T<�����8U��xH�]�k�8� V�����<����"��Z8�?Ӂ�s-/% �H�u��� ��h�Kf�K?���?{SA�L�"P* *RY��T�%|R�O׿#��U J��z=E��"�#�~�ܫ2���[�k����l��9L0���G�/�;���֞V�q���x;)[����	��JWoWx,���q$�K_xx��7|�x" ���������chj�F42��]�������p�1���,�Ns����3��Ap�1�&G"">��Ǒ�����X8��6��d�����x�Q;S�ڛ����np;ꄠģ�	EXabk�Ѵւe���{"����T�P�g���Mh'|J��>��a^���� :H�E�,cPG	�C
��w�1v
�w'!ӥl=���on�܇��s��r��q]�'�мͶ�Ӊ��f�}sc�P�N����D�BoNcF<�� ��[w��Oc��]��v|nb���+�;P��E7��["����S�DJ�x�Fޙ�0�^��IB������U��(S���0�5>��xU��s�o������V���0+��y!�"
��9(�kD��0Z��ѿ���kװt�6.^����0�����)��O��w������)T5�#-��9���2�U֢����������G�	�c
D�vx�v�05�����m��DW�0��s�����$"-�I�J)@Nj>���PZ���|Զ���sgѶҏ��F�V>��Bh;Ӄ�?����x�/?�ݿ|��~{l''�^������O��9�����{p<u����>^�t��Sj�ԍ�	�fR�'J  �^P�x@U�!�
2��P)§Z'	�2�җ���"4n������Y�!�����DZ[��	Z^��\�X�I��Z_��� �1���(A� �A�6��u��7�ߙ�4w����y��om��.��{'��׏z)Ym��n�C���VE��&A�ImMÑ�8���P\��c�+�E�t+��{i,<���V��hؗF* ��z��,G�eaJ�J�,��</���dM(�� J)����L�g5�P�߰԰�"l�B�JC`R�����\*R �#� G%�G�8SN��0�G��2^� ԉ�1G�p�G���W�2ר6F�a=�:�4��e���*K�q[2LYJ��.����W!�4b��K�WaN�Pn�e��z�o�.�l��D�1�},:x4���x.�4�["��E�=ɘ+ƽv�H��*Irɜ���*��g=�H�xm �JI�<,�rJ��jk��{@)�:	���<��w(^O	��썂�x=��
�=��D>߁�ߥ����-�R��A�+���5P*^P�N�C���?T�6�}d���h����hg{`;��o(���y%c�a��9�0ec>��A�x�Z�$ϔB@u�h=�"�-��f]��W�6�M�0i�?�x���0cݑ���V#t�Q'��߆Э[���xAǳ��y����L1<�����S���.A�z�����e��%p��e
B�TYO�n|�9J�mg:�D�p��W�s]U���B��5#j����ٗWB�ku���O�W��g��_~��N#�<6��0�u�e�l���67YG�Q���"dM�!}�
�(ZhB5��� :Ϗ���x �z~Hy@����FBh�~Ԟ�W!��<�x��W�)!��Z^J�����Q}�`�>W�W��Q�mJ8�$��$BoӾ��+c8�\�Z����6�Bp %�H����^ S�����W�^��>^E�W��"`�]�yCe*55%�A�t��L��O���W ���o�g�
8/�����V'ӭH���֋=���h����j���p�6�,K�!t�=�
�J�N��3��U)��q^7�P���so^��.s�&J�P�/\�C�a�gKW3��l�aKup%pz����Σ�@Be`h ��q<<��G��A,C����H?���H�Eو	=�0//�xy"6��<��io/'{x8����v֒8�憴ٌa�`���P�g&#$�xN��Ζ�i�`K�����Y3s5�L���M��� �(D��|*�P4PB���5��*��.���MC�/��C��r}j3
?�$�|�dl�wT<����0��y{V�wx,�O�t�]Ʉ;��4�B�&7��(���/��Na���q��Ѿ;���v4�y�<ӇA���7�0r�zkS�h�8B��po����y���X�=����9t��Kƀ���΃M�����T~��:��2���>5�9���$yB�,K�@� �:E�=ݘQ�_x]yA��,�ְ�b�y=��㻸������Ɲ_��ƣmd�g�-���>.GlE*�[�P9؎�)lݸ��O����[ϟbpi����G����'�w�̭�@uS'���	�U��iEAi�22�8w�
����Ɲ;��Q�pW��1��4>�֮n��u�`EE5HN�Cb\.br������|h�@�rQ_R����7�����U��,FJAu�J�:?��7q��y�/�֟�ǅ�]�ş_%��V��V>!����٨^>��b� �Pݽ����?@�	�+�ٮ>��:���#�k>4�DJ���� �o�P�j<��PY�D�=u(�c��g�]�TKաl��[]�:;�����;7�֕����c]B]`�C�Jjo+=xFy�P4^��ƀ^B���.��#��R�]��N*�ݷ6qr���p>R�c��#��8֒�#��)iK%���X!���{>š�/���LˢƁFÕ��$/҆��jCq-����PO3���Y���J�F�@��s�t�i�T�)]�5Ga�5 ���P��b�����8?P�_�f����Qc�p̅�P.!T#������:Q� ԙ �=_��Mp#�* 嵔P\I<dҘ�<�Fn�L0di���Y'�ڶ$��R������ޚ�g¤/�F�f�a U��A���&$u%(��ڨ��!��x�h�+}B#�%}��h��!4��QJ!TB&U!m�J.��) *�Ò�T>:[x/	���o���$��4��7��SO�|
|��4+��)	�^��@_�P�A �R�QՁ�ԋg�wT T��j=�/!TƄ꼢�C����
7��H ��� t�z5�����_S�g�1��t(�Y0Ʉ���P�^G>O����3�ϝ��>�Pc�	T@T�T Ԡ)��;��^�j�5ߟ��Qj��F�4!�T;"w[���*c@]&�^�'�w����,��t̄7�;�d,褌��Ǳ�*/�!b�Y�9�)��� ��w�� ��6��RxTG˔dJ_�9]Nͅ���ה���\y�
���O��vo� ��}J�7l�Ù�8�J�#e|���2
!�Șk@�t-�x���:TJ��SC�4���#h��8/���&�4_F��Ԝ�U�Ywq�p֋�S�Γͪ�>K(<ݦ��gBgå��s]��(�)a���i��?��v���%Ʉ
 $ u *^MO]��n:��4��W�r�|_<��2NTM#�E��6�� p�xF�KV�n���IIXn��N��7�7���b�eRy?_���i��Bp�sE}�<�2����M��-,?����;��Ͽ��9��^��	l��
�J����=���u���C|G��&tO��k����T�!['8�����nޮ�;櫀S`38�N�Pߣ���󄻏�
��	�Dxt0b�#����%B�r���T���ą� �h �CrH(�{҆�����5\m��Fu�ʅ���� ?wd��#7'A����bGG;8<�����~����$�4�0Tðl\-����`$�'!����-���H�����M��_$j s����`�$�ꦷ ��Me�]�@��)c=ey��O��]|	�b�O�3�)����I�{��K�}�@���ԍU���D�v/�W�����gM t� :��Pɢ+*��2t���|�$��a�$�Nߐ,�н�N�P��oīu�p'��@��3?��3�\��/��?�����5�x��S���u��f����Ta��a =��}��z���+��t��|+�n�����̧��%,WiT�F��T.e��L�}<�P�>�]]�W�:�K<�<h��
N}yw��.��c��O>�������V	�q��p�s�U���Q�U���4Mvcro3�kh@iG+��;�>:���!T��e�7���U��z+'� �����97�����E~i	�{{�����Z�GKW�*7��[�;s�3��FKK�2�����(UL2�	�I9T&�RsP�]���TW����yMH��D�X=�=�w��<��_���?_\���\���"g��M�|DP�����sB�S^��S��X^��'���@�%�M�=������
By��		��� �p��U���JJ7��2����dD�&QR�D5 ۟�8�3���*o�K %�r]\W*bi��0I�A�6��,v�9�س���M�_�D�z#����rf 3�V1ve37�1pr��e�:� �9��"�5�H#��<���Q��II�p����@<������gf#�?�Ȃ�L\}�>��Mܻ��MBpG<*�;����M�	�LCPk�;�ږ���8�W��%�	np���,�9!p��KI��JV�oAhI8l�5I��Y�Jf\B�yQ�Z'u����!�S	O%�U2)�z?5�)�R՜���Cou�CBp�L�#���
D��T�d.S5_`�f~NjZ*�^CT"��h�#|"B��3\ ��|��)uֆ⺌�P�( �Jy͕!p�.}��H��YS	��� 5!|ʸO* j�NC�9^�ޚ��Z�gk�|f��Щ�4�I�x��2ⶔ,��F�dɒkH����)c\�E�u�h�~)}ʠ�j#�Q��Q0: �rB<�B�	�^)@����������yH�쨚u��4lӀ�
�Վ�P[�x6%���㩓�Ǔ�$�zJ�Z�`��f�rnM�t ���I�3���z-|�0өП!԰�|��}G
n)�[��:�4_���H��~G��RJ��NÄ9�v\�e(Д2NT�2���PJ�Q-��'T_ �R^��)���Jڦ~����>�:�㚠�N���)t�A�!}�9��`��A�`(��������>�@��_�ܵR�P���U�{ܸ�� j��yO�9rg?�^��M�0ܵj��"��"�W��0�>���މ�N�Oסl�G���\���F����H1v�Q|}����+A�l5�MW�K�L/��Z����`	���~+��P�v�/m�Nr�;ʿ7��?9�S�)���O��/����5DK���cpi��[g*�Z�a���X������B
�3a�i��kkP�����]W�f�*��� "��L�*m�8�ƋC*W�ު�	�{MJU��:�[��nԟ�B�9�"%ˍ�5M	��T�y=[�~y���1BIB!Y'P�Bp��L�n
p��S�S��H�u
p������6�%�\X٧xAbe:ɖ+���y	���%���k�U�nbقΛ�*	�
��`�%�ʸ��ԛ�kƀʴ W~�$ᐄ�
x�dY`T2��}�G�<�uY��il���2ns�=�P�$m�q������\��7��"�,�y������9�Ď�d�-��!�p𷇍��-��noWx���hP B#���aA8�w/W�Lݼ\p$����	@iE!*��������hd!9)�٨�.GNz2���!������X���������no;�'���Ow�!G}P^����T������$ۮ=���ioG�g��:'Xq�Z[K�K^K��u=ꌐ�`ĕ�!�=	���X#7����cP�˘Ї�$0�?]��{�xj��
a�ך`*�r%c�AP2�S��d�@Gn�?�Ѓ �J�m�	qDgd&�7�y^
@w�c���ooa��2zΌ�i�5k-
@�������_��q�	w�I�k%���[���Ul����O��)X��p�3��J��� @�R��w^��}@I��;�w5���l�A�B'���W^�&��S�@>(�� #c<u�=�x����P������ޝ�,����8��)���y���ǯ������W��˻���Ddy4���X�����#u�^���Wg�93���$��'2��H.,���.n=z���a$#�a��Gw7��������3�.`fy�C�8qz�^ƍ�n��ӿų�_<�=�HO�GpP,"Ò����$Ą' <(�>G������' �$U�ܛ���W���O��/���|�˿��?���?`��\��2�����K�C��%L?#T>�~<�-��]�Ct�����@7?�x@Ub"I1�RQM���( -#��Nd#v�h&��z@_y?��~@hd���'�9U���dL"�0�C�( H��գt�E�h�����I�]f�*cF��ӓ�0�J;���-U�lM�oى<E���z���yv�����C�HҺyn	(����++x�����������*q�������7��w�0#�F��1=YoO�Gq�\`� ��p�D��(��Qp,&�R����*�eQ�baSF�$��\���1�dE��W�sV�%7fP��c���YpU�!	��B�A��b jTJ"��t j\� T<�����0�:�L�"_�	�Ӕ�iVt�1j�#���@|G
�I � ��w@�9p(/T* �Cc0� ��>u jD 5R�>	��OQ��5�S�]1�qcl��<��V<�����K�!!T�7�?�ɘ��H���i(+�Mh1��-�~�}4��]�nQ§���N4���/����Lÿ%B+Bc�Q�~�Af+�o�q�T�s�@(KI0���O5u�.�V���K2D��<�����4�L��-��z%_��ȿ�t �Z�|�xO��P-p�K����D��w��ο7 �B����P�t � T��pܗ�PB��Ս��Ҵ�������e�P���������H����"m�����I_���(�m� :L �}�gK �}��V�	Ս����HB5�C�v>�mP�?�9��͟e6��K}�����_,��h&��_&!r�̇��'%I�B%�{B�h!L.U#���f��滪!�H��S�YkU��z�aO0�*D �Г��ܙ��,�v���7N�ƩW�~g£+G��*F�V/�?>�O��C|�X���ȦT8��¡)6�]�򞋂S[
B&�;S���
��uH'��@�W��zn�W�	b�$DMgf��󒀈u����1�5���3�	����<ق��f�: � �A���:�M�"��Dx�7SmK��j���Z����B:��
��s�6�:��N�waS�2W�Ћ����xgu Z��|5 *��؎��#�5,~L`���k ��)^O�y��T6\�WT$ *���T��'�������Y��g����pR��hQr��tɆċ'PY�%!Rc?ߚQ@:��*��N!Wr$��[���;��=N�v�����_o7�>� ���������� ����>���c��-���$�GzQQA{,;Y�HM�Es}�k����� $DD"56yii����������77x�������q#y%y�HK���icmkk�;����.N�up��-����m`cE ���9,�M`jm+s��z"4㸚� �=MkM��1�ͧ��{��@]�<XD/��@9F{wL�m>�iY�c)����mH�!|j�݊�������7�c� Ti��, :~{��3^$��* ]�����+�9;���nT�6�j�	-��i��� :��ޞRc?5�@g1/᷼�[ܟ��Ե	��h��L�" ��i����������+8���� ��h',+ ݾG*�;���?�j TA'�C`E$	���%����q���O	��йg��9/�C^�3����yö?�ś���/�__�7����O��?Ý�C�B�3��>����8����L��vb|ws�	
��b��)LcrU��hĵw���ӧx���>U5���������������7����ǿ�9�:��p��<���=�+o����	�u�```�u���@��_�<�"�x�S�������$�䠵���������s|�O�����G����y�o�$��)������ǛX~_�X�u[&|��<����Y����}� ��V��b�}��O��M�>�W:+a�\?��;�v0r������ID�[�;	��~�p��r�1! Z���"�h�g��7O]�@!�2o��0Z��-v��eg9���o�ﭠ��ʶQ��I>T�ӬR���1���U�����
BS�R�`BOt��n�X�-��	����hB\;�p�{���PB����8��eBKL6����OU���^	��Xx�ǩ���%Q
@m�	�O�"ea(3�0k�������2VԚuR�eʪ$�\!T�peQ5݊B)���R j�@�l�^�j!����n52�ad���P���^��+��) (PYp%�w0_��·�d���(��Ӄ �1Qw���f;y=��� Ն���p<MT¡4���+��H��&��%F�4�	�Cߑ�p�� ��B�iҀ>$�A�q�o1��.�i؋���I�{���CJ�����>*/TExTstj2��0�	�R��{��멅O�΃������N�"R�wj% �O �'��|�߂ϗ���@"e����VMq�a ��l e��P�id��ʔ{ B�Jxn/u0W���>����mҵW.���&))��]Kgߡ4xP�&�5�����@�	��C��N��|�y9&T��:��J6j�2N�#��O"L���S Ը1�i8�\�BR�^�k�P
��|���.��$8��%��e��9���"5K�B%Bk�Ԉ��*�BFK:W�H�Ŭ� d���E��;ͽ7�=�O7Օ��,8���q��PW�[{<	�MIh\jŝ/����>��s�\_CPu�B	�	
>���ޭ���@y�	���b���jh�T-�7:�N���AL��H�p;���]% "|��,��$D���֞iG5���*e�َ� ZO� T�Pe�ժ�׶r��#0��RJ�R�\�PY���)�F�� ��(�H@���=�YO�N	�������	�j��[	�N���L���t���4,KP	ÕeM�:�>�R�)v��/�L���z
x* %��<W�Y T T����Na���b+\��d륧S4���|���ne�g��3� �����~1�\�\�h+s8y�*�M�����?o���1������3�(/wxr�	��F��	I1���@_'�:[PS]���<�>�z:0�ׅ��T�1a�HKH ��!9&��NO''�'�����c>>���q_Ć* ����7��Q�G����涖��'p::����N.�N[�XZ�Κ�����̬``�G5��;8�����hMF�tV�b��s��L�v2G���%�$�	�Cd����1@W4Dؔ��Ԇ־�OOJ�%a���H<��c�҆������;��z��S/�c��6�@�����=?�zh�R=�Y٩�W�wc�w�0����~�P	� �$DcW�0|aH�ܛd)�!��~|���t�W�	���� �P T�ݾ?��{8�ʘ�iB�����(�@�ai�|j��/����̲$0<'tR����M�`����	\��E<������_�_��o��?���Q>Z�����Nq�o�;+�Q1P���NL�/��݋���۸��[ػy��Kؽ~O������-}�N_�������'�_�_���	�����u�l��ܕX;��������كή~��� .6v��
K����{�)~��_�g?�1~����g�ٟ|�_�����|�Ͽ�ÿ|��?���o.a��s���v>��&_h+/$+�x	~O�g�k�K 4���:�|��P ]z����k��x/����2�ه܆�):��0|o�P�4,�2�~{� ڙBM%�f y(i#P�h2����N�p�%ТE��'����2LK��P�Z��m�d��}}-��P�٨�_98K�^���)�Ɏ��ڨ����4��O�?�;��s~����_��KӨ �D��#�.<���D6�!�=� *����d�HBxo:b�s?\������Ç�L�_M2<*��T�	�-�T�PK.��\�5�p�K�CEl���՚�jEY��4�%A� xZ<E�&��Kcm"�4,�� Ԅ`�}e��<���1
<8-[ba��� ��>�CaZ��p�פ�@���B*�J� %|
�z��
�9Z /§�d�P���4כ^����^1�\.��}�����|Zs�V��0g�4ʁ	۪�P��6_��P* J��`8���Zl��@��NXP:`�������V���	�jC"��	�2^O<��P%�e�S���"tJ�	���5!��q�
<)�ܞ
6��c<U���@|��@��?���`��r��,�?,}�����P�^K��_I�UcE5R ��U *�P�S��E7^����������y,�zy,J��u<�B�x,)}i�J��/󀆹�;�}9�t�z�ZU"0
�h� �҅���s5�	�Z���F|o�rٺ#�-�0m�����R���G�v#�.�!�TV+�Po�G2�d��"�zJF��\���|�|'D�F�
4U���j+�W?�S�j9q��������e� ��wf;	��<{��@��֟C ̀+�ӹ.ne�h^iË_��?�W����kol�_"d
���5V����J�;.����"���6V�܉:�V�h���OۙQ��O���#�:�>\�d��ܦK\yDM���~��\�J ��d�m<'^K�G�N�M���^�k�ZI�C�,�iD�n3*�\A�U�k��: ��.�V��SzV5 z�{*� � ���g� ���)�)I�Z	�:�Tɇ���f�%!"�6^�B�Q�˟�0\���fUa���.u��S���̷j(T3m�N0����I��ا�G8(ՔO$W���S��T"��#*����/��4m�lK�ef��l13333K���m��1f��0V*�pquWuUwW�7��3�|�گ�(�\������+y����{�Zk�-`Zp��mI0��
�Xl���b��Eذy%6o^�-��-�6`��uX�n֭_�ի	���a�F¡�V<m�Y���&�OS3#�;����aa(-�CuU	b�B��h/WG��@SZ�`���۬���
w{;8�Xc��U0�9������7�`-�g�J�r����M밉\QY������oJ��sc,X��-�����t�2,'�.����9�'��-���z�0c�4�,��u�����
��m����ܒ�����Nk�Ped�I:D@,��x<� ���ˤ��D��.|J�[�LOP����h�h�Z��* =�QI��o@��( � G@��?�C�lC�N{rJ ���PN���(8\�Rhٱ*���0\�P5˱:���z��2h��Zm�A����Q��6���;�����q ;�<�����У� U�ԷI�^��h* �^nR�.IXS�
+>Y���dCeg�C�h�S����(A�J-j�
��r�:�o=�.գ� ��k��JX��a\��U|�W���������?}��FJcֻ,�b��0�4�k��������\T�jк�u:܎�����3��G��o�(zwo��ￅO�����:<}�.�A�P�{Q�\��������[P^U���rTV�";�f�v�ŉ#��W��{�`��!��������o�������x��U�~��<ۍ�G#x2��'C��k�Ӎ�[h�L�S��5�붙��4&	��~�G(_��˭�%���Ӎ�x=��Z��'����D���[-|zõ�e *^Pw+�-�{����'գ�^,}ؠ$Bj�����X�K?Ѫ@Ն�AD]��# ���'�&��amqϽ��(��Ҹ4mG>��7l"�����w��nĽ����;�q�d��a��Q�Hs�e��@9m�i+B�y�3a��k�CY[0b������.��倕Q�XN-��#l�b�dɍvĚDw�K�$��r�B>���(O����'tΏ���1/��f����R%"��W��d+�5�>�%��*�MG2��"�����b��S��$�h=�	�m	\�}"-U�yA&XJ`4&��3�6�aKy�@׍�z����`���z�@�hKC4�yީ t.���g�#|�d�A'�s)�|�e��� �.�C�R�
��y�G�[B-!��r�I�ω0:��L�/�L�|F�PD��Q��5����P�(ێ�V�3	��Z�
ӕ�}��>�ӳ.	�,%��E�-�p�1��!��?&�O	�%|j��>��&J%�.��; �8|ά���)����St�N/c]���Y���9��A�6w�����'TyC,��f:*����ER
�j%�3�xM��ߑ<�S�&�h���NL/�,OnO�/���R3�$��yfj%}��T�!TJB�JR$!�9�|�]1�Z����X���	�$S5atq�;�:ba=���8�����H����E�x"�n�	�� �&��&���waۀ5E���)�iD5�D+���ef�q�;jѐ êH�����,O���4/���Ae6q�Յ~X��ՙX���v��/��o��_����\C��^�%8a����wt~�#�����7V��s�un ��cP���h�T�!�1�C�?R�@���1�X�@�P��2��+����>��� @����a�e�@�{�	�ic *%!s̃)P9�������J�!�c���L��ء�L��S T$��6�S�r�x�O��#�G5[��
��8�9�Jt���E�6I>�{� *	682>�%�-�tI:4�W��ؠ����O�$|\�P�>4r��b�Z&���/ �<�L��D�����=T��n�g��ۯ��讞�b��j��AO<��6����:�5+�v�Jl$�>-,L�����`�V��
Fm���h��P�t�bx�1�!p�?/T�8'�.0X��������L`�n-,7oTYqm`�k0\��V��牏F��+�Rvv��z���&?t��Z�G�u����-[	��x��X�K-����X�?��31{�4�ҟ�ً�Ao�4�5�[#����;��M�(�W�]U�.��ʘ��|���8X2��IUC�p�D�p;�t+^O��W����j����/�* ���!ؖ�D��Nl��]���j�u��p�w� �7�-���LU��W��C�(9N�����U)I�ZϷ�� Z��U�$!RС��1H x:�!�賽�E��I�/(t�v��;��ڣ͂{�}7��1p�}��2����%!�|+��m�!�h7+T���t�E\>�J$T��1���z�~�/_ IB�$�7�|�=���O�����V��'x>_P��l��<�� �MH$�����c�V_�C��:�h=�	9W%���`���+z��Rw����=���^��:����տ���x�/����EpQ ��	���vֻ�<����ɋDxA��3�Ր�,�iA+?���h$ �0	��ΎD\^,�JSQ�\��*�v7���M}�((�F��.\�x��T>��S�������R�B��?�o�����]���.��m��G��=	�{�u��;�h�?�>H����ԯ �X�Vqz\�e�d�r�8%$V����U��m���#��1���z���->|V��� ��x�"[�����%������4��>�' �d�-��TA�w��NPzŁ��@ �%�9�:�TB�+m7���~��@�W�CE���BDC�k��2G`%��*2�	C��B�7�"�1F)�EB�ۙ���$��#c$�l��٨�� �i�M��HrG��\�u�uQeNq���z����,�Vv��<����Oc��!�ʂ�g˶|_���$��	.�m����Uʵ��q�XC �!tB�+�,|e���2��mX$��Cm��R`T'��k	=�n�0*�ϙa��P��N�7Ĭ�-���"�������&N`�3�3d��XcL�!�R3	���nv���b�N�P��d	��9��83�Ӕ �n�������q�S(�c��߀Չ�`�{i�����l�N�V�B?���,(Kj���Zm�`��@3,�u�Qa0�KBaP�c8y�7>7�b�� ����I��¼9	�uq0����Z���k��44c����Hk���x��4<S�i�X���,^g�e{�8���\o,���#|�-����Z#��]�9\6�:���*��f�J�XҀ�!�9���e9sl��+����teԏy��E��qo��>�l�JX%5޷/{��`)Ra�/S.�I_�1ϧ��"������i5���i�̊1U�_��"an�&�D=�N��
�}��w�I��$M�~Q�a�F�:��;�S��G�@S ��(.�YÒ�)i��Pw�d��*��$ͨ�:��d���(���y�Q�X��?t���4�'T[N/�3�i%��4���,ه�N��b*B��yUR�9�9W�6%�ie��$�'�\D��,y�ʵ���j߫qo����kf�/(�')���<��K~�g�a53[;v��<w�--,p���,�V!�sR�=*�yg",�S��:["��� I��T��`���@�s�]��ʵ�N�7���*� �X��DakY��c+e^��p,%X.Nr!d\��^꛵"�KiD/�V��cE�#�\Q�]��o]�k�>��7���x?,������~;�0��KqP�[�}����8^%Q�-�BPu�Zӑ����h���D�7��)ðH�m����R;�C���@w�	�qO�t���
��Дu����ꢇ2EX��KAD�v~l���@� �x1���6[���)l�e�@%��)0)����"�vf*�@e;�*�	���T��r|9n%!�*�� ���3"〦#�H	j����n/�ov�~%�vYl]혞���y�Pq� z���T��IBts]T;��r7^��6qF�ji�+I&����C�`*�'UF_�)'|d�.AT["�iw�p\��{�_���kb��l!|nٺ^y?7n\����Ժ�~�f�!�Mahd3KDEG#!1���pvvVrp�'�������F{���A��fe��jYaR��lk	���৴�h+�y^�ka�v,�l���V��M7���K⢄�H�9�cՊ�����ן�ڭ�miDLr""�PTY����^��tt�p�d�]L-Ă���Y0�	���@g�L�!��.���Vk�L�M��_�/�Qs��uީ�W�|����w�y/Ki'|����{K�ʨ��e�q��L|�K-??�L����[��W�b;�V�֠�HZy�G��C�4��$����`�wV#�/-I�h��*c��Y��_��#�(>R���	�TP��=�FM�&��*A![��Nz4���;0�d۟���g����~�QJ t��^�߁�[|8	�M�Zyq��5���C��K���eR��� �G ���lB� (p�9��z�����:B�Y	#��!�4}�	>�	>���V�wx��E���O	�<�
:�I���4�sb¡*���9Q|y'�技� h��ixëB�p�	�xz���EIJ�ܭ��K��
��9�W�����{�B����q��kh<Ҁ��|M1�z%�m������a��,������9~�L��{2_���9���Y^�@|E4��P����<�נ���ŵ�>�;�©����O~������N�#���5~��Op��8��>�l>��w��U��C���.t��䇊�G�Q����3,���cB�$ia��9I�*� �|I*�����?�^�D��*�lU�?�� �Ώ����G=�W�ci���<_�/�א�7A]�p"�ڕ�î����P7��`t{�|z�] ��W��k�7��󂳄�@%;��Ö�jW�{��P�'B�Ù�N��.�/�B\����6'#�6�e�('|�dzl>�"�`� �i�&�Q�!�ƴ�"�=��)�HC6�<66.c�ps��3�]��p�����$nC�ǚpjc�${ T���	��ׂ��(��N��dF�O�Xd��2���!�`�:�=6cM��ƺ� �FQN<�V�Y]a����X�m�E~fXh�E���������.S c��a��H���B7��G�/S
1$���:[0'l3fQ�#0� :�p8��9��Ӹ~^��ƚbn�	t�̱ �:̹��mN	��I�%��R-1'���$�
K���-�����^���ﺐ����Z�����m%����*�X�sl�0�j.f����CL),��|��:�&ؘ������`}`�g¶.&��RB�,���Bl��Z���5�Ì��G��0k�]�<��1͆�	C=L3[�iV�1�v5�ٯ����	��6`��Fm���-Q�[�PK,/�Ǫ���@�h��X�f����*)͘�|0���-R����S��<����h&��*vQoҌ1/�d��Vڱ�{�$Y�d:e9��[P��r��0*���OɄ��)59�h
�T"D� B�K%��Q<�~A�/�K��$�Y��_�_����9'��9��4I3D5��x]c����%(i�<L�tB��� XN� ���e��R���HH��U��I��J�����h���5�����ٟ�
������[��?�L#�N+�:y�y�:�.�/sX'�N��9nJ2����B�p�c�Y.b[�'��v��d������L�co&�#aD7Ebc����b-t�u9���m�.3��yc,L�[UK�D��:��Ѱ����Ժ6Zi�a��=�.��>S	�)�XF�\��j�dN7LpG�p�?8����Ž���Hcy?��C'���z��X�쌅q�X������E½,
>ձlHBdg&rvW��P#�v�!i�@h��2�[)��=@x�!H�"f{�JB$ð�4c�q��ܝO�������0	�"ı��$`FR����ij]ho2��	�l�Ƿ������H T��v%N��iJK��U$�V�S���S��I)�<�ym��������xe:��,^ZY/��Ap�@�h6����F�@�^hh/	�H�ɜ��]+��{�z�W��0*m7��Ύ�6����~�Hx�y��g[%��8A[��HDج�ԁ�+]���QI -�25�m��z{��R���l��������V],]����c��5شus#�	��ϵ��bͺ�,	�7������0�v���l���p�T~A������A!Ahn��XU/o�l�,��ܬdD����V�[��po�CN��`�u���1��p3�n\S�-p��A��7B��ho������"<}�AeMR3�������"��e"!)������9�t�x�2�/&t/���(�-��y�u1k�,�\ �m��tGpF |3��Җ��h��M�=|��I �E��r����g�T�� X�	dN�d͕}J�֫i�s�c\h����kyo�Q'+�F���� �����Y�d*7�`gRzs��(h|o2F��E��Pt�
���Q@,G�Zt\�FוT�Dٞ2�G�0m��v=۩��;^ۍ=������J �1���h;���tZ.�a�T+ �s���F��^J<��i ����ա T ����ɏ��
Vz�
�
���g-A�� *Q	]�H(�$	�J��*�-��K�r���K@�G��]A��7��/�ݿy���gx��ŝ�������yn]E|1C`e��X�	=7c=�u���m#�z�����m�OMq�3��2�
����KEfC14���ęk<ߧ?�/��O�o��������?�?���x��۸xo?�����C8F�����L m�߁�{�h�CI�4�]���If�N�"Y�`s����>�m()�UvA�b�]���8�W�Jޗ�����|�z�Q��pF���8��Ԝ'�r?�~֍%�Jޝ����� �P��/�Bٰ۰a�k����P��)�Pg��ྐ�(� ;��NGj"�z�|�~��� 0b��Q��%!(���`�k�����
T�������!8$v$ �#�݉�b���k ��o�4��Ƶ;Gp��!��]��\l2~�Y%;�"�Me�5����.Z ͖ag���[��+	wB��d"���_cl	�b�M>fX�f��.[��uיa��1:��B�X��]���Li��1��1�s��m���f���
2�|�&�u�7a��Z�t[��k1�kfz��,�U��:�'��R����5��0#�qZ/Ȁ%�� ;�`�)wM0��E��N�/�(Br���"��6���`�v�����T;��(,GU\���X�7%Aӕ�ʮtd�E!���-���P:�z!t,b��J�n�u[��"7Cl�r��偍��Xc�U��^��b%K,&��XcY�6��`C���;bY��G�Aφ`�q!����L�X�h���6l�ֺ[b��9ָY`��9�`���{�a]�C������=�հ8+d �� ̯
��
_̢fW�an9KNO��%���ӳ*E��Λ�JH�'�S�t|^A�tV�+fS3K�4�g�Q/}�B'i�At2��sf�w%}��\�<'HA'�s���Ҡ��q ����
�/��� t��:�C�T�ct���
J�����
B9?�/��p:A/P��$�'��ŋ9I3�3�L�t�)�W�ǜqM��j�-��2�/�)��d�P�M
>�Xټ&��*3������˶f5���l��@u�\�m�b�[K�0����1�v��m(�}i
@E��O(�s}e�KT�I����hXD�B	�֒��>f��"|:����#V�8l��j��Z���\?l,Ċ,O�kR=��]�b�P9���7���/���w�y_'L	�ӽ6A� :�׬��E���QVXg���� �W���zI�'�*	��%t���XƳ�&l�G�3z0������D��(	��WrF����R�ܝ�����p=���@��S��O��XB���]Zo�X�n���C�@��>�Z ���1��Bg�X�-Ӕ�S�Q�@���@��GU!�,���$�P� �&ڣu׻hC�����.���#�}M7$����ue<�V��G��>�<ۮ����|��NԜ!h@k	�'i��,�+�h��NT��J���6x3Jiӗ�4gZQ��!��01����]7+V/��-k	��	�Rn���002���)L�Ladbcz�&�`����pv󅽃��}���_�@8;ɐ+�F|b<��K���++3©#�R⑞�@?8�[���)|���}?M7m��捄OC�l����0$o�4����	�~��Ylٲ�����'��ȱ(��FNAR	���Q(��ŉ����a�E�`���jlP����t1,Y݅z��xt�a�¹�5&�ч��	����_�eŻJ�{s��;PJ{Yy/�%65���@h���\U*%k��P	� �0��'IBTu��ШA��.�|� Z��@s�U�y��(�]���BD�$�>�	}��h!��p5
W���LWH+��V��PZv���2hU+ �� ���;1��.���{	��tH�s���t���'���
�S*w�����v�҉>�
��X?�Y���z@�H%�(�g�)-�*o��!��rj����N�2t���9�j�	�J)�P�V��n�IX�ӃV��� m��}�e�to�����?����k��ï�/��'x������g�{a�5��$�+�@��	��	n����?�VaV���{�'jRѴ��o���.㫿�������?ǟ������>��_��Ï/���q��(���ǁ]�{�#���s�	]wZ���̈́φۭh�ъF�u#������f_���(���^&IBk��9�
D���U�cT�>U\&|(�THt+Z.�) =��1l2
͹:%IDT/���Jr*�&��DP{$�i0�@��	���G�@�4�
�ظ����I�t&�:	��0��c�'$����J\$�(�K��P�!R`R�҇r@i��M���?�ӷ��Z��P�9�)�6�ܿ,���ф"�!Q�Q�	FX](b[c�] �HK����D�93�[O����8|��^0���8��=6�ZÌ��d�����)�ؚ��l7�d@������8G؄[�jI`4��=� b�,7�n�F���b�[�`8m���V�`��f��ۀ-�F0�����6��b�h��²	L����sk�g�,b�d�5�s6�`�7�}#��X��+�6b%�g�e�A�6��`��6�c#��>�[b�	p6Xd�E��X�o }��XO�\O���[���)�1Yn�/	D{s����F<�Ї�g{��\��ǫ���<���~?��<�}����~��U��5��~��2�­��b%�l���;'�!�M�]�/��D�e#�&nټ�U��ނ���<8���z$6W "#��h���k?|���������ǿ�O�|����?������_�����o�_��_�/�����������W޻��P��	V�xc��E��Э	*?��K�]�iuZͬ%�j�1� :���l��3i�� e� T<B4ԧ��av�V�h���(�a/^P����Y8ַo,��d,�R%����ϟֻ9Q3����(5��ϧ�vN/��F����r�����9�{��� �d��:̬�=���m��^���,�[�Щ�q�:�f��)M/�6�At"tN�T���񾯦�`N�3?�9Yӫ	��KO�Î�ʗ@��L�w3B�� �u&�B�����)òzA�:�+��C��+���Cs�=���󋼱����"�Y����.��o�^�#���e8���j�� t�&����h�P[%4� ��2ƵZ�&f5��jQN��Ӿ)n�mH�QI(���"`S� ��0,Oo�֤�ca�օnC�V|����ş|�;o�B�:�s��0��97�:I�����6X��UA�+c�Y��D�'"�-�{h�iBƎR�	�24IRwIB�R�Yb�
@����x:(�˙�+I��
`�0E�^4>/���P9�xSw�!R��N�U�.��:T����������L��N���.$P�<�vJ���Bh<a�e�Z��2v� ��BE�5Ў��J����+
@|^�>/�z�|�6!!TBr_݅�{�ivA3�pHi�JBL��V�'��e��Ӵ�N� �;6��Xb�z:X�U_��V�ش� �i-�`fa
S��eNYp�ƖNX��F�������@��i�Fml���_?�䣴����037AxX0
򲐜M�t �Z!��9�I�ؼW� �n�	%YoM�n���1l,�agcgGDG�����agg���*<|-�]H��CPx4bӐ�S��j�u���ɳ�r�"�c��d���E˖b�rN/��<�:��Q=�ҝ�9�c�Ű�DH�?s�VJ�QI���`S<�2]�{��z���cZrF2沜$�T���>׈r	�%|���T *Yp�/w�h74�ϊ�(���?Z�L�L�]j���L�����)*<�Вc�����Q.?P�����* Z�� ��JBp�c�Q>�������}�ϧxA��?�( �z@��J ���m;���N�K8�C�)ɇ�������߃�;��PI�C�	�h�L��i�q=�z@	���������j�߅O_<^���
ýՁ��\.��lCӝN��:$�ҭNtHG�lǁw��g���Wp����ˇx����'��9����'�ҟ��/��?}����G��?�k�|w�|��_'ǰ��~v7>����.>�o_���������~�?��>���}\|�v]���]�Ix��z�V��[M8�������A�l�ل��aYw����������X/-��d؜J�;�{*�T����P�G��I� �V>+����	�G_�6B���At��A�' *�Y'���,ɩ$)U��l�tD��F�C�;K<�T�Ip$L�)�ta��^Bȟ ��
@'���;����Zy=�TO�H� ��e!.�� �~��@¨��(�E2=���^~�,��W�/|K�P��$�n�7��|Z�m+�ac�eNk`i��#]x��>ܼ�W��DV)�M0'�%�b3���,��1a6&�*��j�̏vQ0�۳Q?\��VQu,
��QT���D��#.#9Eq(,�Gqi<����Mc.F�������|4vU�������l)EU[)
�3Q�Q���
?9����4�4gC�]��a:w5�����U(i�Gzi"�	l񹑈�
ATf0"3�����@�f������L}���|��{�膠�P�5e �&>ɶp�0��3�QKcj�p!����Cx�D><Ӄ:te�\�'W����Q|�p�zr _<=�Ϩ=;�/�n}��I���Q����ۇ˗w�����|�.�;�K_��g���O����q��M�}����=�������C�~�	���'����O��Wx㧟q�3|��o��?�S���o��c���	���W�[�ſQ�B���?s�_Բ���/��U��4�'8a1�W�� �V(��r���[���Zͪ��Z�*�SM@��Y`t����<�3<�b�D���}G��"I��@۞@iG�{<i�$��V��|.'jF��C4]����IIX'!S��L��
�^ �qM��qʔ�p���t*��Wh�^��+˦�^�Ǚ��E�:�ғ;E�j���yBދ�����M�I� T�7I3�</ȝ�)����T����"xj�����͠�'��R�<W)� :���Z�{@�)����`�nO�jY}���Ur1�W����~X@(���P�g�tӜ���]��n�6�] ��O�MWl��	�q0m�V2k�Q���<��&�TU(���aN�E]4��b`U��P�V���"�\��¼"
�!X��%I�X�ꆍi^Xl�����~v>����W��t��X��=7C7^��`N�6̍��>�e�v�T ��(�T�¯V��e���~������<����N�L�Q��i�ù��� ��~j�2�98�@E�L�q"�N�� T�M�SH��EĠ^��S)��*!���}Z�	t��[¨x>>s%�=%QɄ+���~`�Bqcx<��}�qүu
 ��Ah�J �6���	&2N��ɒ�C"�j���j�i�K��xA�U�� ��e��9u�L�O�RC�^�|��C*����T%�4��䃪��*�;��Uk��U����bL�ad�[�6c��f�������>cS3kebWl6���678{������$E��;��nptr����**�s�.��&s�=bc�PZ��ĸ(�8n#�Z#:$I�Q��b@��3�f[9�e+l-��dg[kk�89!$(���Q��j`���0T�ԣ�������M��/m��hd����)y�����ܾ�޾XK�]�|��\N�\H ]@(%�
�.��yfBo�l�1\�H'���;�ɭI��}h�A��J��cQ5�I�9�j�G��rɘK�Z�-��^�-%|
�*�� *}@+O�U�\��s��=J;�X!�y;*�֟��D���������jPrD����;H�Oy@�Q�y�Z��ǩEž
��}�?\�i��c`�����E���t<��У�*w��v��P��Ӎ�,��{���� �:߁n���O��%�N��R�O�Ϫ��l�����dZs����T<���S�ryah�����J��V�]�C�+��K��4��@3�N�|��u<�V�����A��߇]Ϥ��n����{p��p�x�O��ݿ� ?��/���_��P�����9�L������❿~u7����?���!��`��N^kD�+U X��`]�i���ܪF߽z��lD�m~���䚛�x��7�okv�?T"	������9.�|�'��c<Wt�4}�F��$OP��&�jTr�64��i�#�$ �>����!�2� �d�-�8K᱈�BBh�;��	��HI6$��.}?	�/x@,ٰ?�RB�@�����ϱc��d�}�C �/%d>E��%x:}���驖��(��'��і��ea�=�ބP�B?x�n9�p�v�G�;��� ���QVX��q�=я�7���ݸzm7�\v!�0�4�U���|JPS����f���+}C��[�����x��9ܺw�o��}��==��㕋{x�#x��<�w
���ǅS#8y�?����?����sx���x�&=���7N�ҕ#�>ڌ={;p�pFw��o@���z�֠������ $�V�˰��������EYQ2���Q[����N���(�1�Tf��"�A"R�	�)~H#W5碹��v�ȉ4�d#)�
Y��ަX)�+��qs_5�������N|q������ ~zw~��n���7wG��a|~w_=܁���_?مO����{�ٳ�����Ã���[��o?����7��_���͗��W���>ď�>!l~����������1���}���w�ڇ��ï?�o�����������;��w�������5~�׿ß�����ᛟ}����7���=��~����/�_|�>{�����O>|�K��E�aPg>��]�OvAutk����u!����`�n����0��`ZK ���l���h��$��o�t�7��p"��	��M��oǁ�.�c��B�������p9Y2��d��(5̊��J�BL�OB�T�>E��蹦�,�/�N��� tf���B�zAC��k�j"x�kr�h5|���[Y6�҃ ��P��|)��>��o��l�o�fTI�$�o�fP��s@g򹟬5�O�k�|wDө"ߥ�@��7wL:J��YN`%|�,��Y��M�X6�E�a*���b�BD���l�t�&��rǼL75D�|~��xc!�W�S2�Kح/țpcO��IQ๕�1l�Yk,,��5��jX����&ƕ���M�U�����TG�Râ�Jq�~�-�$:aI��gz�(; ���`Hcz��.����x�O���O�������zP���� ]��~��D�r�U�Sa(�Y�j�ӓ�ʓ�Q�v�>����L����Z���&�(P��NyD�Q�٪���JX������GsԼ��j=��MB�8xj���A �PY6�^�)�i��r���=P�<�V��|�\������)y�$S Ն�J����@	��� m�����2!��Rm�B�D��S@l��k]萱?o���Β��H ���a�tS�7Q��cYn�Zs��vy+��D��G%�y�)ڊGVC_c�7�������h)6[n���x;M`jnB����A!!���Aph8��ݸ|�l=aj�'_ls򁃫����������4����ή�z��{�������Q�(.�#�F@m�JŅ�!���[�`ih��[`�� �F&�O8l��5A4,$�HII���?l�h�SPUӄ��R�x���/a1)�M�Anq5�+j�SX���\i	:�QXV	G',\��W����%�p܅���:�#�.X���3��d&�n[��4o��"�"5��ۃh��ɺg=��*bGK$a3�՗����{N� ���^�je����1t�
eG+�z�s�h�����P	��,BL� �4�����]�Fh�S���/EUs��|~�/�y9P��=e�9�<�#
@��ȓ��A��N�T�o	�G	K��O��֐���M*E�Dh��v�=��I�d�>����v<@�Yq����@�>����Vz�u���x?���������D���)^PP)�Z)C�L��a�@5����t~�(GƼ���+|(���B���!��f4�jE�m�Jf�v�R�Z�}�u��u����:����A�� ?����w���c{_ߍo�S:��!|g�u�����`��v{�7P��V��k�h�VCؕ��w��Z�ݩ��"�s�j���(]�o�B�o3�d���K�^��I���D�Tu� �0\����xP���$�~�%}>%s�H���r�����Yu�
էkP}����I ���'c�Jvd�H����Ng,�ٰ����V�E�� h�'�r���G��l��`I	X
h:���v�P-p*`KR$�;ԃ��) Jp�+
@@�x:�L���'R���H�L T$�aUQ��� �6�QJ�\$ [��������)�"��ç4�q�X�Q���ׂ{���޽#8u��e0�X� 8�zyI@�)a���`��a��@�"��ڔ�������sc.����c���^�{�_=���O���'����x��aܽ�w	���:��{o?�����3�p��N���۱��rt������E�h)Rӭ�h��B�F���LTf'�:7u��/JGe^J��QU���$TĠ47���(ˏGqn,�8ƢJ�F��ĩ�8��y��F&������<\�'G����&�y�	�i�g{�#�)����������0~L}}w_���W,E������>�я��ߛW���\�_���޹�o�yo�y�|�:����x��.�?��>}�|�	~@��ӏ�����?�?����S�ٟ�?�ɧx���x��-<zvO�~H�|��?x�g<Ɠ���O��Ï����Y>�#�{�������C��~�O��(?އe��XV�5-��J�k]_
�8�h��*��B %�@�P�	��iLϢ��y��pDe�Wx`b�@�A4�`0�T	��UJ(�0N�H�M���3�N���I �4��TH)%p5b*y�H@LBQ�^ 1����s	�E��
*�(��/�&�r�x;'i�M�f��t�����>QRG���R�~U}�<a�`=� . :Y�|��s�K�xO.�u��*���,�R3�ߪ�:VR3y�T�_	)�p�J�9�%!��Ǽ��3�9�g��b9����Z>��u,'i:׉f�q;�3�A�<�}:5�V�>� *�U#��c��,�gP�+�[�E�|7C��.�,�*���&���^X��%~�a;�O]Z�UaXC-����t7l�
�N�fścq��
� 5k�Q!�[�B��FM�`\	CM��TD��U"���k��P\���L<���0)	��t,����Dg�Jr�Q�=`���z�}�����}���v�(�	������y2��S'��b� 〺UDõ$�mx�����*h��V��W 4y�d�-F
!4ig�M<����Aݞ�����gR$���S��HȮ$'n;�T$�0�!��>��)^P��o׏�屵 Z� 4K�ݎ��
� C@�����f�yH�=��+�{%�v<�P��|UJ�R�
�ƨk�N�ud!�X%j�v��F�*>��H�2I4C �����f��M��~4_�Q�����n4_�B���h���Ӯ ��ԡ�SC�^Bn��rxn��t������`n�V+�`�|�0\��ƫ��d=��	�f���T�O''£+��������
D�$`����R�v􁙍;���O_�_d�/DBb&||����������_~��	��
Q��� ol�4���#�hY����6&�SK�����.�0ᴅ�%"#���c�'����v�(��GCs���G��3� ��̂J���iA��	�%Uh����G��ۏ���88aͦMX�~=�X�Ka�"}�_�G���i��?K6��!�ay�(Abs"*�נ�Z7�a�,U+P¨��s2B%�ZJ�G��/��fT�^��M�\%!:+I��TІ�-��~�� ڎZB��hJ��"}� Q�Ɉ�NG��{_�O��EϢ�UQIJT��c5h8עru^�B��JT�@��zLx8���#�:�h#�J6�t��ʂ������t��>!H �j?:	�]
B���S�cPV���Y�Uy?k/7�D�����|�����9�h�b@�rՄAUR�:Bi-��;h�ۈ���ǻ�h�݌�j'aU�u�����v�o6��F3�;	�|��vq�0{��<W+��F=��C+�L U���JM7Ѩ�z�V)��x͕W�;��) ��A(d���Y �e�) �|Ac�) P�t;Y꼓��O�5~�ΰ~�W�J<��}@��L�_m@E�9�sߓ��(�k�Y��2�\Y |�X�ʔ���|+���,Oʙp*�pe�l�I�(��;�<�
�[��R�J�T
F?������B\}$�_U�ZZ�(6��5q��$ �:���b��А&�
�z�x����[���`X%:`��V8D;�sw#>;� ��v�G��w3�l��X';�8�	���0�v�i����LS�`k�ԺT8������N�_�};*�k��7cρ6��cׁV�9?���q��Νą3#8~�gN�����ێ���>ڂ������(�wlo��p#��18P���Z��i��Y����P{���P�MYj���P���jBiQ�3�e*
�9F�CqNʊbQVB��JBskv���@	b���`��8Ct��Z_.�m/�C-�����wN���K=��6���N|�`'���?y�߼���#�����3��#�6��E@�=��;�%�/�A��Z>�ҋ����6��u��.�?܆�'�q��>\>�g/��W�����p��~
'n����q��U��'o��#�N���p���zr�q�ۧp��B��t���Q캴#M�`�֢���;��~�>��'��O�Ư��7�����S#X����X���=�Xݕ�%4D�4A�]�G��nS�9����1��D UIV& �H `� � ��w��
.'���Y��Mo��e�dL+��dp�C��P(���1 U}&E�T�Iz)����q��������x�I�(P9lN������5L�~Rڡf>�p^���m�PmH���/ :��)ĐgK�5n#���S� ��A�' K��>��j���z+��hLe��<]����@��L��l�h�R�E�n* �Y�wB�'�iĜ�`�i�� ���� n��L��L<���zf5����|�R��B�:s*�W�$��0�W��,(���@����y.L�2aԚ���(
<?5$��b/,�s��*�R���Zw&��[P��1�פ>
F5� � T���k�ۆ�1��iu4��VY�=slL�cs*���m����pl�w�Y�\�Bм��>~��>}w�^Gϡ>D�c�Ӻ���M���j���̱4�V�ຖG��8,���MCwo
��!y _��I�v�>�j,PBh���WI�D��������8�J)�)˾��o��F��"���N�8�d��1B�G�y=��:@��Q�w�\��8t�>��T *I�$W T<�rы * -�ũ
@siI�!P	���T�I6\�$���+�h�ک����k!�6�M UYp	��:T2"�Ӧ�2K�zE�o��k�^�΢3���r��G����M����po���u�b���6��C��OGgGx���� ?�@D�& 7��2->��v���l\����n���E�@_.�
�L��w j��7�8{�������<�������v���0��|����������ؒp�7O��*yx�"2*���0������<���������DE�"&%�Z�:�V7��C"�����W1��0:���V�X�z�Z	��K1�*a��P�Y��p:tŴ��Fx%�"(Ǐ�b���Ps�Qկ��h�T�}"���*�%W�s@��ͩ�2 �V}@w?>��W��ڞh	��� ڕ���	 J�V *P�R�ud����C[I���P-'1��� �c���?�15��ۮ T�~6�!0�a��Cy@���J�.>�����������aeu�i�� T�5H�J����T�%�xH��K9��oh��o*�@ʗ�z�Ѻ��h�E ���Vo 6�M@�6��N+�ﶡ�^;�գ�V=?|��M���&? 7Dmj��`���6<nԢ�z�ՠ��Y���.k	�2�i�f%㴊Ь�\+���_�~�S�I�61��+�v�U5>����B_���9|N��򉒏X-�-���,m��J��[���X�O͙Z�^h�f�P^_��z����/q��kG@U��.RM�c�T.
�t�%�OY|J�M �"�y�+�;��6��O��tPi0B��.�B��݊׳4L�gDe$�+"_����<dt�a�t���x��"��#�:U��Vư�f�c��'��,���k�*�M��J��]���n�>�}�����ه��$�P�D{�����kF�6��@	���0�BRe<�\?�[7�����W��������6Y��H,
G6���-ń�̼`�&�#� �E(�L@�X���<4�V�e���"�4E���h�DCG4ͅ�l�CYm6
*�P\��*�Wj2QQ�N�L��:U�(�Fv���ܐ���T�{���MYnr�}����\?�$9��q)��NGn�5v5%���R�.��%x��o��燯t��C���(>#�~�p7�y�?~u7��<$���7\�������~y}_��ל��� �m�'W��6�_�S�з�h?>߉kGq��S����X�$"%?�5YH��D��;?��S˓V��g(>ّ��o��v�e�L�l`��H��6�b��X�k�����i�%�f�uߊ�~fXh�g:o��۟����S|�����_�m'�	��R��0��s��
d�sa�4��G���Nc��D�{����$�ʴ ��O�o��7J�@xQ��F;��I���S�`���	lN�36����8\~���I4>8�3�N���%�L	����)A�e�񿏦I��$��C�,u�I���&p9Y���3�rf�>g�n�P-PjAR���P��|�z�tΩ�T�]��O��<g�/*��s̮���_�ޘ5.ցh&�t,H�y/g7)��e�ٔ�ӹ�d=߾�����-�P�j�j���4�b.˹|��4+���9���+��M��o����T`isV�'`amt+1��K뢱�&��°�Z)�u���mO5쇊��4�Yޘ�℅�NR��bf��:�~���HJ�O	���P�U!��mP��8X@�5��y�����Wa���Ȫ*�l\Z�a�6cK��G;as�Ǚ!�;҇7?y��>߸����d���Љ�!��) Չ���03��Yp���T� hTW6�wW�`-�F���p@�a�/�q���$�	����¥�WPN��4�;!=����l'���]�Bg��+�L�Ɣ�:�̷ҿ��Fy���� ��� h
�-����}���3b��4�D���)��ȸLƍT z�CŢ͂ۦ�R�S��
�	��l�:o�U�@h�˸���}E����}/c~�Ҟ/��UG��p)"����~��\�ś`��0��
S+c������.N��Gl</-iYHNIW�YRZ�Ҳj�'g��'ޡI�ɄwHBc���r�����D$����N�hln��[�������7!00U�UHMJ������H�����������6洑-a����q���~����ߣ��I)وK���ͦ��z��h����'�|"x=��L�D*��shU����sc'����Ю���������	I0��ƚ-[�P�q�B�J�P]�,����Y��a��>l����ڕQ-1�<��t�l�=/�D ���=�P-�q)}<�55�JP�Frܾ׎��� j��?ю�#-*������4����T��dJ.9�Q Zv�Ň*Pt��\'《T �z�K<�/P�* �z�Mg[��S�v��
���{/�^���f3�YQ]��������jWP�|J�[�O�7�[	�* ��M� ��M �"��*/�.�F\�C�,#�U_�y��<7xLJ��Z��q���]��z�i�&�-��T0ڌƛ|n֢����`�t�A:�_�J M���>�ohx.� Zu��	�n��2܌�6����X}I�NJ�C�I��X�0��#&�۞��p,/P�N�8�* [&�YÏ�d��Ũ��5\懑�o�G��Z'?�]h��ʏa�R�+���R*��z�jQ�� ��)�'�F�1�	Exm"�h���%x����@X�V���2%Y.�U��h�d>%P��
|���!�
c�J-���I����C�3��ttuR�S�ؘ�X.����"���"䅕�p�8�#`�Hp�V^T�\x�z�O����>���n����W�7Z�����øu� dМ�H8��s�5,2S�`��2�&y0�r�A�L�ac�ԪD�����S=ر���X��x#"��)npMp�K��l����2��r�yJ��ah�p[8��r�t s:ԁ˝��g������*���m�-`�l�l_s8{��e#l���y�
�n@��r��A�kj�B{a�3Q���4OD�Q��m�ӑo�98?��;�q�?���h_�i�[�����A|vg?���=؃/��_;��x�,�쭓���������N|zm?�ԏR�q���g�F������� >�����~r��_��;�:�����.Dh������i�n3?s���6ESI�ؔ���0���EN �s��6bf9��4�U���]�b��Ls_�i�1+�3�1�w�$:bi��%�`������uv|�>�����_�?��?���#�G �s��%^��4�[�X~�}.�b}o
�I�򂊁�$a���D#]B�4Te�T���b�,(�H  $L�
y$XN��͜A����S�f��&�����&��x���ʽ N�K-|j�Se���P��%�M�@ڴ���"|�� (�p�$������W�S�Ǚ 9�L��dIȭ��8|�b��S�h���B跡��<���c�~�3����W��}0� *���(��8潤��� 9�)XIy2	��\ s&At�s�f�zٮ�PI� m�ܶ��7&��芚á��L�.
�۪q]�r.�sYkVu$b�&�[ba8�����X�vlqu8V5�A������¤=k��*�2��YX����v��d����\����(��`�@����,PiKE���T\Ps���A0.���e�h�s�6`�#T�ȴ4۪baU�M�.X�m�m1>>��<��_���>z���Z��wP��󢬵a�]~���p,-��\���:�{�!�hK
R�K�G�N�^��0\Bh2!T��67��-@�hG�s�g�X�τ�yc�?��E�osb��� *�He�O��
���4��3�f<|Ӷ�2sg�J�"�#��B�^-lN��)t�T�� ��.^Z�4�x�������=�*͹z�VC;��z�Ɔ˴��tk=�*�V2�v�$D�������6�ҡ ���Y#�I���l3��4��?J�:�W"�ϓO�/�}�h�|,߼�������f025���<�<D�KAv.�)+�y�ͩ��L����!q���LG@d�����,l�a���08@�|C��փ���#..�l�����&d�����v�V�
EX@0\��Ùǰ2����5�,�q��,h���sWx��/�u�`�zcTִ��>Gw�n����CHt&|B���Ϡ$g���	5��h��G��.t@5�mP�^C#a:[x=K֯�⵫����L�Kt�30k�4�[3[�6#0��/����ڗ��/9��6�w ��u��&�����?�}�JW7�h�|��/�,�2h��f��h{*b:h�J\���O5��x-�%� ����L��*4�!ۜ���D����H"���y��/�:x�P�S T �:�|P�E��v@�|6+��"|v4� m�Ѫ��5rZ ���$�YG� P��� ��	�rΉ�[.�Py}�}�����X<f5���YÏ�t�f��o�����H m��ȏD�5W��1�$K�D-?��{Q���\�$���!��t��7�Q~��>�W�0@��o�§�Nh$���x�	��"P�p+��
h����Ys��D��r��i���9V��R ��H��w�kS��i�l�_���|&��j�K�t����]�B;�̗������A�������֫~��v�<�FZ�x(FJ_
b�b��%!�!
@�k,	����pB�QRF�Q���DTuKQ�ZN � d�c���eZ��gD9aVJ6�4�éH�`!4��rH1�+���CTU�Ҡ�`%YTNE��w2:��]��uCx?~�~j g�lO��ԕP���4_h�Kp��.ܿ��Ad��4�u�5��]a)�
|f��(�ƔI�+̒aj�����v ����Ihw/�Lw�r�c��#��)ΰIv��`i�hB#�M.���B�l�c��:lr߈u���~V;�g����e+6�)��Z筪��f�͞&��a��N���r)�-�fӅ�wZ�`d�9��(�[3p���Jp}�wv4�Ξ6Bf5�S=�d0�F3P�h�=ͱ�B����"ܥ�o/��Exx��N6�݋����(����<9�_�y?}v_?:��?:�o��'L��{��Ʃ�y�o�����{�!�������"A��>�2��@�v��c�S�]j��|�����hn+B\n<S�����`X�G��)��*�EMl��.�:�۰�`�8��S\���
�7����>x�|o����n��ʂ��$��9���Z��A��>��'���~�O�5�����87l-	�z�O tz)���{�f�zc�&�Fp(��Pn�Q�HC��D)�7�����W�� T%}[����aE�MIH�]�:���"lVO�ɐ���� �\.p�]�&��8̼@e��� �����_��`hr���t*�|�^ Oo^���;��e�j	����S(�5��لϗ���s�|��J��!�Ʒלj/>�<n�1��C��v
x�M|
x�m�Ǽ� �k�փ)�9� 9� )�i����Щ t�xH'@��#�t(��H�Q���Ԫ-�8�V-h��H,$�.n��nm(5E������.K��X���"�O��%l����ZX�ee�Xƶeۀu��XS����*wi���*��9��j���,xv3aB 5���qm$��-2ei�ySM8�*B`@ 5,	�AQ 6lMkb�К��dذ]3+��1�2�pXRS}���&����߉�o��G���7����j��1����EZA7�z���#m`��-���* n�!
���� Z���l�� ��HM$�*>�/��b$�)A�N%�)@��B�'3u_�R�<�OS�R$`*@*`:.�d�幏T"��u�r��)B��b��A��aT�lD��r�� ���X�T�Y��j�g�ͥQ.����*��h�Ϩa鋚��J���NmGڇ������J"ɝR���hߵ��WI�BiK
������M��v��Z�Z�r�W��v���M
@KN�!�x��"�3)�Xa�6��:��04�S3���-������ 5ngRJ�s�T���K-@i���(�h@@L�����[w��N����������ܾIi�	�GW7��k ��Q����;C� ?X������!!Ox��!"(�!p�����L���e��M���ꋈ�q.�����.\���~�5�4m�MBTB��zں�������l�U[?;�ڷ}�{�=���T6��� �%��pt$�oĒ��h�JB�b�-���KfCg��Z1����'�"L��#���E��P�b��˝�E�� �d@���P�G�?@Ǉai�>��)�\A��&h��`ga8�i��HA��T�$k��sv�%�5(��W�E��0,����x�|v��;���<���a�<Ŏǻ���.�<ޭ̀�<�v������g���w�� ��m�M�����)�o{����Z��3��e9p�üH%�t��3t�����z�M% �SBq�Pp��H��H�Fn�x���C����:�Fy�d]����~��ZV�H��	E�;Q�P�o��@�V�VA�6TU��R����儰
§H���*��^o�A�zO����#Ў:9��UG�|EWDͨ#��^#x_����x
+`(������U�WBjųI���s��w~������xŃ�i��Z���E��� �xY�/�xX�z	�*��9�7Vo��z�4<����Bhe�JVa�S<�R>�F��9h�7^l#l�>S2=q��J'گp����}�u>78/������R{���-�<��h��Z����7M�?M �*�$YdK|	�-�EX�V��ߪL8� �?����.�G����Qal�ä����� D�sY�C8�hjle$btK���(�jh!�)AXA0Rj�ٔ���|t�!^�s�\�����+!Џ\s6؆�V��q�����\�{���+F��F�.��P�4gX@-��aJP�e��4��&H$�;?���.!�v�EJ�?#�a�m�<aM`2��R^T«M����`e����u���e=V@��`C�16�RfX�i��^�X�k���Xh�5A�X�g�՞�R���X����݀�K4UG��H.�,�u���J<=P�G��po{�>N�;7�C���\�u�Pc�]uq8ٓ��ù��������h&�/��#�q��^��7�����g]�?��U���,w���xr������Z<<X�j��|tm?}�,>{�8>����{Wz��x�J޻�c_j�;Z�V��o�Sxt��֢�+�%��"<:�>:6%¦1	VI0��6���mm<VgxA'r��aE�gzB�u����,*�C�At^�?��à��w^���^��n��o��~���+����||���R�U�4����BY	��*?m�4B笆 趄C�9�2���%tI�����3	u�d��w*�5k�d^e����_��k�>��\*t�@�Zϥ ��%��u�5UH���5L���ATP����F�d��w��;�3�\�}M�q�:ƔP:��n$�U4GT����5ҷ���b5����AOT��J�-��S�9�߸��Y��*o,�%D�f�]1���G%�q{].��z�j̯���:�'$�'$Ϋ��jnc !T<�|����k���}nSA1s9?��3	�3	�3�L��v�����eJ���9��)�Ix��<��������+�E�c����,j�Ţ6�Y����B��W�k"��,f�xb�&k�	�XӒ�u��|�c��1��C��m���0,�?Jq�E%����ӗ�|�W2!4���aM�k�>;K`ߙ�mm�h$xօ����\惭����?6��u�w=�A<�YE(Lʂa�s��0���e�6G��&�m����{�苷p���7b��,�3��Hk�*��zA�Xn�l_�h�
j_�&"�� � �ƶ!� &�nF���,!���d����&�!}_R��5�;^��)"fS�F$��^�RG�2DJ)����#����Dݙv��܎��`��N4r���+�1r� ���d���H��@��5T���U(9$�A�Qv�E�	��k<�x�d:����k�3x���T��*�ؠ#2&hEU�t�$�sPr���{�|��7�h�IvT�H;�vR��5���Y�.�ݠ�}M�wv���{�Y�gT�V����\�E�m ��p]�l˲�훨�x��/�-&��X�y�mX�M�kabf�m۬ako�m���占�`xz� 95�eH��AZf�����Ņ+�Q�܋��l�y�@���p�AlJ.�{��}�O��	�K*�����<�ֶn�z�����^^�qs���#\l����7�/���sC�_8"�^��>g�������>�!���e"6!	���JL�g�����!Q��BV~#bK����TBq!J4-�s��wAK��w�C��>t􏠡���ٍ�Fx�W�n�
��X�e-�X����Cw�\�,!�.����a�k��� D��"�&�|�{��n��~���;���QF�M�U��-I����!�Q-�nv*A�+e�Yy>�gjPv���|�~7v��@�w[P�K���|��}�#�&�e#_��<E�|;4g�|�J�V�P%#�@��峢�;�9�i�s�F�����'t���J�t�B_݉��*�V��i�܅v>�]�	���|B������@%�m�^Rzϙz�}� �t�d-�S#�AY�J�or�{��ׁ�{=h�M ����� �I�ϧQ�:V���YC Ԉ.I�V��Y#a���N T��p^V�D	�6�$�SA(�F�ËZ�#�ɐ$�}'�C�*D<��w���z|;N�򚫄.�/��BX=o|�9B%?2� �A��:9���P�!T�~��ʋ��M��%�^�sI"���ߊ �k`pU �R�B�P���k��qV�>v=5FKI��wm)���k"�
�*�/)�v��*e�'��Z�v	��� 6\lWY��_i��O`T��#Hu�{y�yZy�f�0M��:h����Z�z�x~�{�a� ��v`�'���t^O/�j\��RQ�Eܗ�p[6�!�>- ���+�S
g�A� �FB�J	�E����}gLy�h�Gxr>�6i��j>�0 y-�(��AVC22�_I(D%��<?�&@	�~<�E��·�4�U=5x��:�~�.�Ene,ܹޙ�h��3�v@M�Fy�0�v��4G�$��Č�$�r�~�٫���8yq���p���U�=�>&9>0���a��=a���OX���,�[��	�FX�+��!�["��5�k�n����cY 4tև�bS�5������l��ixd�ء�*{��qqw9���ݝ��Bp�Ԗ�C9x�=7{8ߝ�#u	�'𺬞�X���+
�6���sqm$�w����<:�������F� ~xw/~x?>{t�|���s
>_=ڊ;�p��yw����U������ ����?����!�||
�!�^��G7����n����>�o>Eo��ƙF<=U�;���oG&��S�7l�UQ0���aE4�XJR��t���U � �K�<�� *Y-���IB����-��McS�ϝ��
�Pt��>���5������?����`� M���\�=��ji��P��	��s�hn��!Tr��ǟ@F8!8h=k�7	��&H��((U�`�R�) ��ĳ8Y�Ǚ$�g��i�s	@NN�3]4���\���<�߅�?^
l�:�����F������~/h��g��S�o��N�R��r\sD�q͝$��Yc:� �[�y�С����+�����
�q���,��@����C7ߕ���A��K����K+��L�eu�X�g|Q}��:�~�G0�[�9|��:�0�3Z�����H��T��a&X�jz�fR3�3�3[B1����6h� m����8,�ǒ1�\����~�Z(j�t#�!�.i�Va��Zb��)
��#Tv�E��X���M�VM��EB�<�K���p��2�����A� ���+*��q���m�g���0kJ�;�ɉ�UǮd8v'DcaP�CB�i}0,���`=j|�����0�2���\����e�0��,*Ca[ۢ X�{"�2'o��_���|�ARE*�:o�B�^�愙C'���a~�	��Z* � -$���k�a��B�^���Z����#�NWY`S�*���]E*7Y twRؙ�ʑ��i�����T�]��=�(�!\z�G�y�F�C覆o���'Gq����so?��6��C6����ߥ���G`�;�-`�	��7�5�1IH��^�O��Ny�#�(��-��C�=�����R�2�G�eB��ʐ2�P�E��hܨ@h����T5��v��Nh��N Pډ����Rm�V�k-W%��W�W�/�.� *@�z�]���,����mձ>��䀞��1�h?�ٶJF������/�z��0����6�m������+|}����p�%� -+9�
>��k1�� �^�����TK'>[��0���G@4RrJ�WR�]���ҍ;hl����=�v�

KaO��vsG�7��	�Pg�NMks;��5,,�y]ΰ�v���3,�l9���xd��"5=!a�v�G��~����W�"8"��y���&V )�6ga+r��PQ�N�<@D��~�:�֞a��®�G���Q�9r��%0t݆Uf���d#��_��k�`�2=�,��y�fc�*]��/�Q�����@zO:�^iG�>���HDq��#�\1�6�v�>��:�P*Q-�R��(�C>�:]�������{�se;��Lt�py�E�UH��Ets
��Ӑ�+ Z��sm�=�s@����@ˏIf]2�QB.�sm�i{�܇�������`����!��@��!�j!t�:|o��E�m>K��7|{� :�����%�v<@e��~���F�� Z�>�� as�t��픔�k�O �A �Ӂ��<��^�]h&�6�Z��FB����T!���.��|�]�Q���MB�������P�M��:�Q=o��o8�c^P��U��(� ���-[	�c$%�Z��J\��1/�$�Q�\�|�`uM�P���MjZ�5�c����:I_�q�V@I�|=��eݵf�d�a�N<��oS����%|Y�P,�U�"V��m p6��4Qr}�||LP�V�^�ɴԑ\�\s����[T�c�s;�z�KI+�0��l%�* �����N�0ʲV~$�����{�q����dZx�F~P���5МѨ��\��!N� %��!����Jy �Ѓ�-�._� 6���Z�q[�Wp.A�
��F(a4�0! JE@��%c JE�#F T��@*enk*��ذTE"�pMp�)Ch�67 �����!��x���'����� R�lo�$��<�E���v��z�O!�"��p!t���P¨$2��0�q��t'�$9`���$\�w?��>��-;߇��`�EZ�2�N�1�E(������5�{Ê��I�#6��`��1�B�����ln��!�X�k���\o�u���g�@+8Y!4��Ah���Ѯ,�٧�kG��ho5��Vwn����`.>:\���8_mKBW�+�<7����f�b�p�)����psg��)���,�����^ħ�O?�H�<����g;qk����C	OO4����M�~|~g��3������C������c���(>�ڃ���=6����6A�-B��g��߻���q�PR�So£�qKA ֗�`#�qM,;��S��g>t!��tg�+t�]1��ɔ�[�|�ts|	�4������ZGx��׎������~��7~�>
F�1ك�	źV�]q���%á��y�4��� �G �����!4����O@"t��&��J����z'��xY����+c�&{3���/��ˤ��N�w<�4�i%뾫�}!�w�=�T�zQ3�@���'H~�x_�qM��� :���II9wL�9��P=�BB�
_,/���"/,�wy)���
=���k�}��е��Y2�j�aV��p�S�R�5��P��uaX����XX�E��ŒH���$��)�5u:��CXp�?�HM�-ɹ�MIB���B���̤f>g���1�H���.��Ҟ,��'Z����TxL��T?P}��H�$�.k%�>>����/�q����:�e�!d��,z�O�eiU(Ua�L��e]-(��2.[L`�����${L��Ă4~B�ԝ
��t8t&8��=
�Us$lZ�`�� 5���Ɵ���Vf8a]���`��7�l���P;�c��x�����?��?������,rX}C�#��@#�1?��l��X�(��9�:�� ו��v��2����Hܑ������� �;�4��4�g6���}��j^�v��� 탓�7�u��T������ z���������d4{j��[���l�6�۲���>b�ۯ�b��Xl4K�F��P�7���M���b!�Ƕ({D�Y���(<(�#>	�����? �W�e�q-U0*�&��1 �#	;���/W���/P��͐���+�ڹ���L�2܊P�c�z���Z/�2��T U��r��;����I����X�^��Xf�K6.�����[���Iy?흜ww/x��!!)��W���Vnߍ�ѽ�i�@uC:FQ�ڏ��������Ĥ#1�1I���MJGAi�ݾ�+�� >>�N������I�$�::�����]`o� K�m�j`��[L��26��=����N.n���Abr
�����(|�����o���n�%�' !�y���}J�DIeJ���4va���8q�:F�#���-�8|�v<�C'Ϣcx�)1Xi�	kͶ`=˥k�@��,��e:*w��ep�#�!�.��	(?�A��!��m*�P�mzq�U���Ra���y�PIJ5��0,��4H��[��~a uG;� ��;��֛� 4�5E���Py�6�x�	�S�dí?C8R���VС�����v5����}�G�v��h�s �@��`֟l$��`���1��+}�إ� ����t"���h�:�B��9<�C'k1�u��;��� v<�C��t��B�����F0��e�t�Rֵ�:��v�S����������4HqZ�3��[wAʱ�O�+�����i�_�:�r��PEI�<�c�*����7��P�A���F��PA.׋gP W^�s^�lf)�)�&�	ї�T)P-��	�Z@�B�d	4
@j���5�<[�*��.��cj�%����6~�D��0I�#�~���r�<��C�f�}z�����������R\��_����_� �8�*/�@�H~�y�S����l�z�t3�@���l�V�_7��ѷ�§g���n~�x}��&��1�=W���hOR�I�!�� Z⁀"7B�L�h����h��O<�s��O�$��ChH���З�L��bB���#����iIFA'�_����&��;����� ���P�%�zB@�*Ba���W6t�(i+ǅ������ە�)Ɔ����b��#��X�����<�	�W��W��w��ɳ���Y��TGXb[�#�r�a��0��U J��{�<��O�%��(�k�-���\�m�~f��k��s��)V��b���x���e3\�.>�	�y!8�S���j����[��wT�.A�NK�wd�?r��p��^B�@�#J	��[��~�4��.�PI8��g�T�����޾r<����r<:V�g��}������On �>���x��������<=ڈ��P>;݀�����������	 C@�����i|~�0>�����_\��{���ΩF�s�	�m�;���M�)!�������y� Gwf���et�/���|n6�9�P�dҔ�Uy��Kv�>��TW襺`^�3��P����W����,���"z�h�'�bE��v�������_�?��?�;��r5X焵|W7E+�R�)�Q��X����'���T�CSz@��9��a.&f�}y5�P���՗J�C������&j.�W�&��'K���&k*�Ra��:ISm�_%9�TP��l;��Mu��4U=H��$tN�8��C�q�:뿕��BT���	�>X[�G��IY('V�Q����mu��[c
�Q#刧q�D�H�YC��
���(F@_��=TǞL�6�aKM�ՆC�&:!��3/�P�o��J ����>J�U��4�j6�u�S�ng<g�G`vG��C��c� ]�� tQg���<�^S�w� ]����|��$$�W�jB��*��5��S⃅�eu�X�	��,!x/��r������� �'��>u��,��G/���an�6��ö=�I0'�ׇc[[�<�&��0��0~��E����T���M<�@�����ް+�e�<r��� �o��.�=���,�[�^[�0�
z�N�%��b�7��@�� Z�m�x@����y�+�:��d�X�P&����>���a��P���(?D�:L{�H�N��>���Qt��C�.�:s�Ԑ���p��=�����	6�o \.���9�Y3��M�lj��|:���%�u�h�\�_77��"=�D�9��'��Il�r��i� �k���Y��]%�aS�4s�,+V�м����2��u@ �;Q��o[��M���:SC�Q�lbۉ��
ա��"�l���@��H��)61ױ���CJ0��� y� �����:t�l�bػ�����w��+����"�eFV.��PU�H ݃�������	o'	�=(���;w�c�j�F��]��K�0G��; م%8w�*v�=���0�Hm8��������s ������%-abb��{�[������pt��HH���!�F�������W 7<R�~�8���;�!鈊/�O`*��x�H��sWӆ�N���{�܅Ԝ"�4w�ąKؾ� �>���c��>���a��:l0ۊ�k�B�>t��`�r]�ҟ	����V�� �-qM	(��!}wh3���I����$|V�-�x_'K2!�>���U8� (�M��
@i��hñ.4��VZ��YE�o�@4m��,�G���^��Pu��r���_��
�zn���n?��h� }<��h>����=mn�~4�k:ӌ������o��r/zT�N����>ע�`�SC�hCp�	���q}�x<%w��9x�#\��fN>ۅ�o�šg;q�����o��~���(�Y��<�v`����tv=!@?ځӔLo(}W����A���yx.���7��2ᖠ�y�ݷ�w���!����J�w�!^:��D W��ҥv�Hn�ƇC����vߔq�x�k���OP&l]�zt[������O�����v0�M�(�xvzM�C
�w��V/:Y_�⩽$��c�!��uܷ��l��@�l�)�Po�B�O$���@)�'L6�AIv�v�K�q��u҃~�y��w��>��j����}��,yoeZ��]mG��^��D/����긍|��e=��1ZYO}��~�{7몓�Bʞl,��d�����d�Nՠ�Bzy{�x<n��̏k��*T���%{�ї�P6����/tE@!?.n���
*�z��T�L�
����PBh4����~�K?D&�	�1�KC\����.�낐L�H��VӲ<"?!پb���p·�B
L���/ۛ �o�2��-���M�_9� ���](�$`[�6���k��B�� h!2�[3\`�䈭�H*O��+���ۗ���qt� 8�6a�
@-�<aF P�l�g� I%��z���E�/L9����*��=���� +��b��6�[a��<�a�c� ���Bq�-������Z<�^�G��xؗ���ɸ֐�Wj�����g��+�e9a��!�v��N���i���Ǳ������th,��c�xL����N��͋����Q��/_���M���\-&|j��H^;ڌ''���ý��^��޾�����Wv��+;��(^?;��#�8ޜ�;#x�H-�>ވ�N4���x�d#��G��3<����xr���������7;��QB�7�"���&�#��2[�㰶$���ϔ�\�C�M��(�b�3�@���.���yX���0��e����3;p�gx�����o���o�E�H��e��5�1��� i\.m��J�/+h�,�W	S�Zh��W�1s1G�� 0̬!�)��P�!�dϡx�XN�������T �2M�*_��^�q�����)���g4���M��_S��e�^Ë ��l;����e��d����H�D�T�fL���������%5�XQ�����rl��ј�ЖD��#���TL{!"�s�V���j�Q��e{ڠ�G�{'�t��p*����p�� yw="G*�ә����Ʋ�@�[ׇA�!T���?´�{@C�TOBi)	�U^RJB�>��9{>gwF* ��e�@�@��Z�N� �/h;�I""J�Z(���Bq��s<Y.��\^��	]��|x�%���X�M��R�#J(կ���$�k���"oB�7�e�@'��򼰄�8����8k��[aC)!� �ԛ�m�	�n��5�Ǫ5�e��`���#a�sl��	��	�[�|�.�[���)
d��	�� t���7�����q��!�7`��,�܂E�PJ7��M0�k��:�����G�Mh�8�B�9{�hԖ��@9JUA#��k�h=ׅ�㴋�*�-e;���^���X�����5�R�e�7X�����at�6)=B�����]6���+�@��˛��+�`�}�!\�ڰ��/��MzXi��Wc��rz�;���i�,B��Z� �Q���
B48EٻKUYx���a
�[�h�d��P ����[���8W����TP�gi�J�'	�U"p���g�U�K�I�y���-J�M��AH�r���f%�QkV���!�Apuu%�9��?��a
E|RrJPR�A���GO_��?�
��C~9a.�
�.=~���w�
�s*�	��8�d!+��Ih���ko��ΞA��y���W�������_OG�;��1?6�@-`j�My?-,��:9����ChTL,�BB`nm���A�����J̄��)YU��d�'W <&��CXL6��xR�Q�Љ#�.c��#(���;���=ãjX�[O����W���MV&�di�U[��Y[D�\�gO3����s�|��y#�-	�I�r�н
@�x�$W��VѾU�&K��4U2"J�%q�� ���tӅf�6��Yd@���>�ȦD$+h9�hU���� U��7�5�P/}@
��Jx{�Ky@��� ��$D���[C�&t�8����i	���'��:��w<�$! � h���t��~���3�C�s��	'�g^ۍS�γ�V:��A}���S#8HH>�by������G^�Gx=�s����O���p��8�� �<݇=���2a�b;�X��E��Cuc����7䶇�8���Ǿ�{���k�Z?���{���o����Z����A��NFna��5zo�>ڃ�<��j�]��^����fBj;��އ#���w�c��jB��7���`/�_�O���~z�0�u�<D�ދ�G�p��8��!n����Ϗq�nv���w��&�v����[�,�oF�A/�x�u��=��8��~5���=|w7����0�w�z�`'��!��0�]�;��~����ay�<ۇ]�O#�X��+�c��v�wൽ��}�����^ȴ��փ�3�8�D��>3��5h����g��1����|�w�!g�Fs�՗�Ț �y#�ċ�� �� h`�+s�
a�L�T��|8��r:�
�qW
��x�p6��H6�Ql�E���R��Oj�sZ�c� 5�@���[��,������`���~�__��2]�twl�7�e�3�����ݳ8{z;r*b`�k|7�� c�� ��MY��D�1Nq�i�6d�e������[����I�B��1�6I0%�e>	��\/��i^�9ZS^�LK�NoIt�j�R��Xj���i	��m0#���n���r2��Q���yx�H���6�w��q�37ړp�)�K�����e�V��Q?�QE�9��φ͂i3Y���`����������Ց\<8X�GG�i��ǃ�����n�����\�W�ģc�����s��Z<;щo^?���{�˯������Gg������w��Q>w��V�Qi���x����Xoo'��Ιv�K�s�M�?=ZC %)č}�8N@noKEZm,|eL��Hl�æ�H�5%cku4I��TW覺@O�~Rs�P ��C#o������s�O�oz���;c��)|�ۯ��O������QO#|}�6�iCp>�iT�7G`qk�IX`_"�wŨ0DI@$��܆`��fՉe���(C\xb�$�!�M�(҂�<ƥ�a2��E*#�زY<6���z9���H������I�Jcp�}4�ƥM�3)����%�5]�s�����Ӌ�7z����E��~~��$ɶ3'I���R��}���:�:6�S�^�T]�l�R���W�M����_�	t��ZX�O�
���@l�	V6���ȉ��CJO12�i�wW#�[�|�����U�6vu���0�����h�މ�]h�Ճֽ}h�ߏ�c#h;���Җ9����y�0:C��.�u�¸1+k°�1�Z��#���.�򝐰�� :�"y_��S�uH;�0�+
s8-�3��uFc~�� :�"P�\��2���͢[��
B�*�*ḒW�hYX�ŵ�XJ0\Z�k�%|a�&:��1
�P	�]X�}�[�9X�6a�$5Ku��XK�K���������e�/�#���}��F����R������R�������Y���mf���q�'��d2�p2���k��n����w�w��{����]���^O���Fؾ��&õ'qR	p��N�v���Hlb{��N�Z�m�[	g����o�4���m�k�{���NcxK��e��6a���))	��7c!K�c�	��^�x@�(;܄���(=\G���[Մ�4|�O4��`�Ҟ��0���m�6��Ym�
s��Ŭ31s�Ә��)̢�,-���k,�d-�r�b�\G�\���,��I�`��/[m���,�x�%��[c���s[�p;h$��3�;V�
�-�G�˕j����@�
ŝO*����i���*;ـL�л�@%J�:%��,�>Bv� qo6�d#y.�OU��a�~?Y�� �^���f 5�߶��o����&�&=�2�SyAY�8�NIDDIH�T�$!R�z��=�pK��R�X�})l��#0�!!A���F@P(b������J�7�����m��GS� J�y�M](�jFZ~%��q�w��� ����Z����W��{�W�FuC+&Μ�W��]4�-?� �c���Mp B��2T ���6��am㤼�;��.^��
P����:}B�ñ�z;:���~���b��?������R��%gV�?Ą�#�Bt�2:qg.�Fc��^T7����EU�س���B}_'<�i[�;b��6,Y��V/!�Zb΢9��x.�V[�/�yYH�HG��t�P����h�-/�M�j����%��y�n%vK���H��7��T]��iS *a�U�������d��*��d&:Q��^%!�kOGl[*2�Pr����>%���Zh��J�[1Q�g�RM��x�3��5�ܨ������I {~�# ��S *I��y#����C�_�E����|�����7�}��}��ݤ�׺p�?ܙ�#���.h=X�V>dU�I(l3��#��v����(�mq���4�/��^�:r�Qԓ���Ԏ�l %��(��B�@��c��������#��d��s�f�����7D������Љ�=�ԇQ��l:�7��/��3m����˽�J��y�h|]���#�}��v��߽G�yv?��x��I:O���xNT��r�D�*4��!l5���W�V{~@΅m�g���~n?ˑ��sw���Ʈ;��1��σ�>C|i�?��48��,e�͛��\+��1�v��Wz0.�MȖe�l��Gkh�֢�l+��c	�\��o�j/Fo~�x٧i��G��@��w������9ߎ��h>V������q��9���,~��Z���\Jc=�?E����ICNW2r	)�CYJ��(�C�|�d�h,ţ�(�]��Ĳs6���.%hʸ΂ B!��q;�(fx�/"f���(�¥V$���O@�~�I�z=���DFv�v�1E��b�
��P�ϣ��1���tF˄Ó����E�r���GP�?�ő*	� ���/R�*��q��y�=wzT���݂m:����`K�/�`6`�ex�:?Xe�uO೔�+���wo�,�c���~I���	�s�0�%�۳xl6d�c#���������`�S2 �6ƺcY�6,�ل-�6���g�#��"���j#Ύ���������r���-9�[����|���|ѓ��~��,?��;x&���Z>C�ߦ{o2#�td�bo�������%x�X-�K����~|��S����>'����i=��0x�dj�{���?�U�篾�7���\�?��k��Ͼ�o�wo�=�k���J�-��)�{,���\��ƮR�-��Sx�B�����g���F�|�ϟ��=�|����@���ל���d�7$��5�����0�D29��]���4�V��[�b�
�5��R�~>5����8wԜ�?�
�����[������h��u�Mc<v�W�b1��e��J���a,!�4��a-IX$�Js$A�`Bx�x�@_ a������r
|��Ȳ �$��fO�,�#��"�H	/ܦ��Jٮ>�m
���D�����O�Q"�ϣ� jJ���1	�	�=��f�6?����$�CP�<�'��h&�y�}R3;?-���/z~�4]���Y�5e;�,�(��u^c�F�L�%��X�I`�`�x<%�jC4��ܟ�@�{
�ܖ�������hCρ�={��]Ëￎ�-|��?ď~�S��w���������������{o���[8{��^=��'0v��^;����ï��~���ӯ���ϣ�30i�m�5-|��-��Z	z���g� 9_�	ٕgE`S��{c1��ꏃ%���q���|ɱ�-xL��OK§%�s~a��95Ԋ0<�� \�y�yuZ�w�s!%�� *I�@�7������܇��T�}IHDh\�>nQA�}���E�2ݓ'�����L/�t�B{�
�J�G�q쌃�͉�iӬ��-6�O��>uKY�@��?���¶BG��$W��%�ύ���c��t w^���cCX��<�a�	������a��36a�q'�A�r=܊��I ��W Z��5'ڑ��q�ccg<ª5pI��֨mX�s��`斧1{�L<�~f�ys��n�s	as�<X����2���e�h9�s�|,]aIYq�c-�>!	���r�m�쐾N�ߴ (m�](!(�h������S�@T�}
�JH�����DJ���ej���ؑ,5�J�H�#�u�������ƀ��C�j�>�G�>4��VКk��"`Lz@%�������2�L�mH&�ݯ��W)�
��d��:%.��[����xEkN�"�3vW�߾ kv�&�y����OOo	�9�-*G{7�Ρ]hn��ȞC8�zG�"����D��ΉI�1��m�8x��+�aH���+���_�����W�il���q��E�e���?Y�Y(��Gl������Q!�~�>
@��&�o]�����~��F[QoP�ᑑX�q�*������?������Sbt�\�V� 3��9�Hϭ�"eJ���c�x�>��U *�o�io��űs��[��ܝЧ'@����kvl��+yoɼ��a�x��u�&�"�?�d�����Π�� Zo�l����x��TzӬ)�'%�P	��q���@	�'*�t�	��ۏ�kch>Ջ�ݓ �@ -"|�#�;y�KQv���z!���PI:$ Zt���ʸ\z�5b���j>R���0�xA�U�]�ӰL�2�gǕ.t��$D#��� t�
��j�*S����C��:�����ùg�p��������g|������ξK���a���VxEn����,�ؤ��~:;��|��l�i�`�RK�Qӓ�f�5�2nKFF��er�M��T�$����H��!���d-�4��T}>�0��H�W�e?*:'q4S�c�\�'xD@�mV �*t�mNDR��|1�*5H��#�9I�(���pv��0��t���˦�˶��}�B2��ϔ�?R��ߝ�G�e���Xd��(e�&?ZNoNB*��X�KR],2Zd=A]N�
UeLY�j+�`!�*$������j�CՔ#Iu&$���V)�����=� :'�R�W���I�8���mj	9�]2�ʺ���G$���`�����"�[�"�{hy-��[���gw��zO9Z�ԣ�X�`�V�\R��zg��"��F�4���4�<#��<�d�-�P,Ʌ��{�T����<^��4�z©��� ^Q�Q���K 52��OP�}R����<�/��Χ
�;�DA[���P����$�����g�<��mex��u���m\��u�y�M������h;�mԖ� ��6��Ö�׽X��P�����/�wϽtZy@��W 4��y�3��6�zB}���ǚ\����zɂȎ]�'�H"
~�mlc���Tv\�`;�yn�_�5Lz'���O��K|�|��1�~��F�q�'��q�F��4���fM�z4G�`�6�ߨ!�����n	�%O�w�,T��q�6	'r��p}8w�q?8TL�,�s'���n�w{>z�*~��5|��8^�h��e��ɳG[���Q|��}������ڙ���7���k|��W��cxp��ǋ���39dRC7cwS".����Xn�8z�x;�����Kx�X;?�	w�7��:\�_�s��0ؑ�����Vj@pU�Rٚ��i!��s��,3ybuj l�6ձXU������9�x���l���Dа���lv��Zq��g�_|���_��＋�}�+�* �6����e��Xޓ�i �p���.fu�i�)�3	`m7�)JBU͞D3T���`6aQ<^OJ�R��i�P�\B��)�'�*^OiG���Tc��
���Ǥ�j
�~^��OIy����i:?)���iz��'��H��tz���w��`+�9��y��� *�iN�y|��Ϻ����ڊH;�p�1!�)�V��(�4Ҍ���7��W��u��?�������/��_��RS����c��?��O��?�'~���#���}�m\��ϟĮc�q�@{��Q��*.�� _���G�=X�]�X������a>3��X2��E}	*Z@ T�p?Pj@��+b��.S¨� ,�(��ꉇ%�A��xA'=�� T��� Kʪɠ��RJ�\	ǕyB%1��:�h�^��.k�15�P��6�B�2t�@h^��.a�� ��	���A��8T�0B�[_2v�����ض���vێj-���i�VD�����p�d�f��cs:�>{G��q�w�u�~�6\L>X�s�7an�vXE�bi��
��1�69a�k�EZ��'�ԙ�̑R�E�8��@숷���e?3�π��<̳���;��r�\��<��.�ⵋ�D�K���Êƽ�".Oj�b,R�<v�ǚ/b��%fYP���\������{'l�a� 4�{j���\�$9{˔�����-��ne��9	��^r��������~����R䣈�  *S�4��F��N�\'l\%d\nF݅F�ۣ�� z�	�JXmz������
x֝��q���H2�
p��o��u\�1���X�]��x=���V�-�2jW���##;�U��kA{�0z�1�����˸��k8{��M\@S��K�O�E`T"�C��4,��Thc3���9|�~����W8r���Kp��5�76!aa���#>�]m<?�M��IC���'�I�u�-A�����(.�"|j��R!�z/�����g�����H�-��7m߄dԣ�� Rˠ��DYM'�+��1��(��}��C�ރBwk� v�ŵ������_����"�0������cŖ�X�Z�WK�[8����Z�eH�OEA�p惫x�����	ڋ�[��[=f��aЩ�CSS�|~ 5{@%�g����� z����=T��%�/Y�E��=^tPգ�L3j�6)��* *^в�5�J�Gk�!����V :5t: �?� ��7^���^�ޛ@e�a��$$��܆�7{p���֍�#��IANybS]��>��!��y�nDx�541v��u�i�C��V�"٦���w�>��zgD蜠5�!����MI�Ci�E9@krC���E�*���U�GP�'�hm&E���a�-��B�v@ h�(;xkm�m?��#��n' �?�t��J�����Am���=|yLp�B=`r�vo�{�\d�,�F�7?��������1.j]Jo=�78#��yD*�,�����<����$_�}�Y^��TR�ĲL�Ad:��e?��Oχe ���BXJ B���d_)�N����p�RJE$ �/`CVA&1���`D$��R�I%�q{�5
le���@�B��鄽� �Ca��>���m�y�BY�-K�l�?���y��8Ԍv��=y0��ұ�2U�ْ�����d�%CEHnH$4G!��$�i, #p
l*��f�,*��,u���R4A,*�[����3�h�5�X	͕�y��}Zl����t�O�/�*�%�8dN���bhh��л�5. 5����5���5\��M}EN�k�lsC�*;�`M�`{q8�z����&u�H�L�����מ�/����*�	�)��<ƭ06lg[v �L���l��VS����	����p�3|`��	��Ή���}�d{���یb~恶�c?co��Ņ�X��4�\{��X:^��Y�h�܊l���0�b��o����>�,�p·,Aw����M4$��$\�������<s�Ϟ�ċ�������������N�eB�ݽ�xpP�	/��G4:���;籫�o�p�Ϗ����7������n��U����8О��c�Mȼy�G�
1ސB M�DO!����H��Ǖ�������J���H{1�k2QT���BJ�\����l$7�"�(["ܱ6�	�b|�=> ���ؑ�uiAX��|ޗeòP�Y��ڦ�����#��M�w�$^���ٿ��|�=��⽠��*�d�D����AY��)�:tD-����B��lU�C8\ئłV��HXp��f�v8)F�I@�1���д��bn���"��E#�;Z-��L>C�{\
�|�ѓ�)?K*�U���4x� #�=���QOw4?C�|4��ǧ�dRӁ�LJ7���|�ҙ�h�g �J(�k8��wV[�������B��:Ԝ\����x��$��"|�����#���������?�O�#a��JUX�q����I=V'����#�����������������S�AC+��F�|��#_���;�෫�;UX�t�$D��3#^N�v�q} ��* �3��
���v��x,�NJ��y-�K$��ٔ�.�+ḄP�V�#-l���#�Z�GaNU�JNdYG���J@T�r-�N�"�Zq+�P�tBD��'ta�/�� �3��x*��k��7���*���y>�q�k��c{<\����'�����J�m�
E�s�w�H�ET]n�}�����{q��y�{�?6h�Lc�yA�0��âH;X�mWc@�Bp]5�(�Rc@c�]}�4xK�M o��S�;6�a]�F�ۀ�˰�e1V�.�r��Xlm�5v+�\�Jˬ0���s��/�kL)�̲�"�ZZ(YR��Լ�B'5G���	���Y`��z�lB]`A{�6O���^�Gƨ$F*T^N�* �)a�. :��H Te��z���iT$���5Oh��"��6O�25T�~�8PɆ�p��@bÕ�"�P��"�T���_lS`Y}�B��q���(�$�N-7^6�Kh��v���q%lY'_�LZDF�!1>���(&|�������6��N����8x����3W�����;t���|�F�!8*a�D����s[��n�׶ ˰��1|��o���I�M|�DF#59z�V��jN;34^���n;k'�$��q&sD�!xph�C"��b�`��'�j���]������͗��1���H�(cY-�O�o�C��4! ̠Ƃ�ִ>���8�k?Z{���n>|^z�����ѣ(���_t$��\����wl���y�.���Y�O�j�l����)@�@>ƞ=��?z�/@��a4_�A=�c9K<�jܧ
����9���ZJ���~� o�Q *!�����`#��K�Й���<d�#{W1
@�?Հ��-�Z2~[z�Zh9�#�P���Q����^܋�/O�;�-���|��W{0���K�Yp���эl���{е� )E��D�v 2z;B�7",d=t�m��މd�LF*�����f 4b�z�q��!P��hA`�r�4Х4=x��Z��vBA18���(���`�#�E�"	�a��!|�bܡ�qalSN0׻�]N@�qE07��zn�o�5��<�=���'����v�xl(���\�uQ���A��r?Ya�al;�0&��8o�p*2����`)�D��0�!Fo�P��� �# r]�����-�N*<!���pD�E 2)a4z���6]:!2%T�˲�Q)a�N$�2����!.+	9z$��P.됐�C<�c3���.)߀��h$p���\�s���VuɅlG$�s?VB�ˍF|>׋b`�e��1�k�DFm
.
�a_��D_�x1��)�AzKrh�KY2P��"T�0�
��N�v�FA�� �f�������L<&��|� ��&����`o������2'!�( /�@��X���4DVa�{[<���58w���>�ƀ�w��/��)�p�q��X�"�Ar{I4�����1�FB��+��կ��_9���u�N�����Y�*W��,�M~0!&6Y^N_8&��-���J�  ��IDAT�I^�N��w��yof� ,���������}-2�n��ǫ�������p�?�;L8��c�a�(	�>�ݢق2�U(؀�H��s����sB�W�q�\�[̀�ay��M�	��\�K���,�?T�g&J���J�L ������C�L_8҈gɴ+��f�za�������|�+'Ǳ��?��K��������g����V�γ'���a|��Sx��AL���<eI��:��R#�����t}/�zp��<�{�N���~�0�]:��w�����8}a?N_>��W�0�w�܇��F�7����uO�WzR±3��/-��B�6-K�"� /�+�iJ�Cy,�n��?�
���o໿������85�k�h��Ij��4r�P�jQ��,B¬�.��m��e㤚©0*�`Q�yeTE ,j�1_M�oU�=5�����*��������_y?նN�J�LiG Tyޞ�Զ�#�%��L�� t��O�N���4��bG3�*�|RO@��])3L���M@w�6��^S�������:��a~�Z"��.�	�j5��1 �4�9Fh�P�U��N��o~����o	�&h�����J�M�7/՟�L��o�_��4�����{���ƿ��7��o��~�]�9w]#h�׋Q>GO"�� B�˰���̔�rB<���j V�N��DX%a�H2,�n1���GQK�.�Rl{ �S��Z6���JPcB@-eh����9B�+J ���لK��y��W<���j=�%���� -�"B�b�M���hqn�JHd��Y�΄Н���D�BđJ�O�+u�I�}g<��DE�2fw�$��(�CI$���a�&\�*�u��B�pr�s�n�m��6��H{��وy��0���%����QӰ���zIB��Ğ\��iU"�{x��6��M;���ƺ�uX�}�c��
,۹�mW`�浰Z��	����`aӂ 9_D�������)��X0�#YQ���	��	��	�f�Y8�y��Xi�An�q��p�w�a�Nt�V�E��2��-Q���5{<)UG��L����u����ʸP�|�8PIL4�+�ό#E(:S�<��m�׫�U��6���S3��P *3>4�N�:ӈ��M���/��GI��T(�S��^�Us�f�Oر+v�B��q�F�@�PTX��l�f����c�q���?v]����9��F��;��=�PXہȸLx���Y�ܲ6�i�@Z^��K��AqE�{����;(����t:r�s�T}X(b	���0�;�@v����Se��E�);��~Ad�H�� 5=A!!p�vGMk5�ݸcJ"�<}�)H�,E|j	£R��J^���Rc@D�3��3���ad�!��Vp%��:�o?�LL�����h��{a����l���+�p�bX.���6V�f���%�ko����w9��o��f?�n����У�����Zq��x��1�p�y��nt�@˩Tj"��1�)�9jh���q�u��}Tw���rBg�D�m'jQq�Zh5���Ò�Hy?�I����{_�$D�&tF�I�|�Mg��}�{Z ���d�g;I�}g��Z'N@;��]Fȉw��dG��A$�S�F�-��	�vH18"�H��q�A�2c�P�#:��)�0D����i�P˱1�J:�3tQr,AT֣��'�M��/?�ƞ7��F��	�Ql'�mF�ݕ�����!PF�	�4�����-�l�q�wr���D��Q�j]�d��A!Q�B���<�H�"t�J�c4A1��M��@2�u��`�C���$�zT���N=���C��"{!26 щ!�N
�.9:�Q	�� ���,�Ll��j ���B�O� &M�J]J��#XF"*)n�������5������0��t�dƤ��ŗ���1�A-�>&EH��S�u\V��2��cY'���~b6a4�`���nP5X�ЧG"&��U�e�iLa�����N �!�'�nFOg��|��������8�N�Gj�	��pD�C�J�-�+27 �s��^���t�ϩeϘ|���Xv�qE|��7�=�l�q����
|�N���3�ڤ��JR��8r������J?�w���2P���O>5&x����26��6�cW��s~$�y?&դ���cx嵋���(vnT!�n1� �\��y;��`�;nsJ����ց�`�^�;���?��K����������g/�+ce�ރ���{cx~4�p� z�<
}�'�����w]���u���$4�B�!�c#�Wc벧`g9I�	����ɦ$\��$�&�b"����ÉR�p�/�jėn��;���gT��#�
@_8ىwn�Ǐ޽���;\���+w�O��"���1�>\��δ��#�xvR/�n&�6��4�P�Q (@׿���4�+��>h-O��}�x��a|��[���^������~�?�����?�3�����;��?�?�������7�������kx�;�v�"�݅��J$Td�P�������υMJ6�i�<+VI>�a+���<8������w?�[_�}�-�^;�pl����N�d��H��.%�."��ǣ��&�Hv��$*�3�07���<1#�ui4NӜ(G�t[0#j#�mx*�	�V�f�����]Kf��E��Q�ߪ�,�i�3�<T������wj�T�#�4���G޻ϡǽ�S�n?%������_�I �����	��~3y�O�in{R�}� � �gi: ��Pj���X����T��OK<�:�����"�?�g�[_ş���	�&5EDN�O0�����������h����<��M�s���_�/��o��ُ�ȾC���Ɉ2�o��׿��� 珡��y}��?;������ځT��OQI��%������4��E#)X<JxK��p,�aI���IP }B�𙌥���iX9��U��X9���)Xڛ�E]|N%Sn�QI�q��:���@If�����2ta]4Hhn!t
@+ÕT�p��dD��C�hB��[Ⱦn�"�sS�1�d����р��ZD���@:���`�b��=v�뱽Z��lw;tg�.|��H�CP��;�׿�&.��s{�{���Z��:b%m�u���
��L�j���@xW�U��O�au24�4��i���-��7	���p���c�;�	̛÷`S�Flڂ-���y�9����UX�����H��Ya�"+X.�$�
\B��#�΃�<�G���[�7T ����������>�����Ԉ��v4��F������S��I/����tJ(.����!k�� ��
Y�ʑJ og4� �"���/~T/Jٛ��~��G��B䟬Tc>[��)IB���!�
@e
�z���̶0�fp��Ђ�ӄ����
�C�,_l��z+�>	��Z2@���c?XO���}iH��6��y-���-�Fdd$m�I�9�m�$p�+o`g��z��;����(o�BM� F�F��A�u��c��;v#��iu�� �e�R�����&|������}���Aff.
r�<�1�����!��`�ٻ���N�n��v�N[DD��K�&*��iP��̜\$$%# 86;�b�������M;l	�Ѵ�S��V�BhbzLI���d T�2�6}25�euh�B��(w��㧱�(�s�A�mq���9]Z
��]�Z t�*,Z��.�Ţ٘�d�m�ٖ��!�K�%h8ہ��A��d@�P��t��φ[=J��	���h��J�g��:4�o����0t{/�N���"A�L�7#k���T54s��*Qr�e�
�����*�ϩy@� Z���eh�>C��|v��#�8������ґ��F0H��;�^���7d+�[<����{��]�[1p�ü!xc��&9݈�3��/ӱ,EF6�zBc4RGi"v��X�\�B 5�^�1�t��F)M4�0�Z����F������^BO�<�h7��G�Ӳ^K����R�'uT�	�g�q�0��N����T��_�#�	�W�p�P�C?3�mG�x#��i�����/��|y��/u��7x?��F�ӍP� ʏ�N�ޟ��7��l�7�~�nк@=�@�K@%\#���q�
@C	����<֝mz�XO�C���A�ć L@uR!֠g�Ueh,-�`KPեi�M'ja���H�Y'���n��O���1R	�TS �D�y|Z�a�)!��$8�T|���l��f�d۱ԘBh��|.RbX�	��N	E(���g^��rP=^��#m�:щV>`M��S���d���s$�-a��:B��p��Z��h�zJ2"�x�?b�Th�����O!Ԑ/� %�x���+S�p�SAQ_��� �VŠ�/y�Z$�%#(Wה@l�8!��7�ҝ�����vW �����
#����[��x����^��h8d��3--Y8ru�{�n�?�}�H)��W�'\	6������G�1/n�Ap%�{�x��nC��F���>��U��n�CT�5��F��f4|��f������Q�v��{�q�!���p��|0��R�5�uZ��[�F��Ȉp�U�[��6��_�3�h�#\1^���&�hN�Ş\��Uv�7���r��雷j�����@_?݄g���p���|�8���޼܏K�Jp��w�=��~�.�h�DO:N�e�|.�f��p..�n��/�k#�n��o��JR�QW����b��ľ>��ų���������L�Wf������W?�&>|�Y|�+/�+o�ĝ�q��~<w�n�=���]��eg]���r�7�#9�Cr��a���tX�ݺ�����(o�3｀�>x��}������ql���r-V��x.j7��X�Ѐ��cRQ	�[�}�O�����g/��(;�<m��byJ�'buj0V�csv$�Kc`�U��2�*��� ,i�aA�Vl��(�����X��i<`A�qF�:R1��h��G���&
3�Ca�g"�h?-���Ow�;O�1��������Nn'H� �>��)=խ�S]O�ۺ�	`�C��)���f�<?u^�{� �)uN��=џ�����'E���������ߦ��L���o������s��|L�Ώ۞f����ӣSz�G�Y��qyv���U��]f����b2�Z�y���(,h�`YU$���)��>�t���k�����3L�KY~\��u��9%	����8vJ��I�_���pީ������_|��Q9ЁΉ��t����_��iXۙ���YX2�F�� |�,	�\_9�=���Be����. �.hL����Oi%at�P
V@	��5W"Ir0����2E�$�gya���J֙%@jQ��r��`I@�O��O��(	�|�U� )�(���1?����X��j~���uĜDW�aߴ�!��p�N�}�	N�q��7��:J���#`[��=�ݒ�`�'��wq��I<��=�3�x_,�Du1NX�eюX�a۰Hc���p�Dyya�/�B���О����Z9�	n1éj��k�?l3ܰ=���w`#!tC�&l�ۈu^��uV8,�����|��D�K��Gӂ`i��r�Y��~J��T+ª%�S�U4o�<���w��0l������dTk&|�"s�L�RB e��y���5�;XE�,G�^��2�6��O��m)c�H�;�e�X��^��"̦�.A�x>a��T��RTH%�Q濿Ս��=JM���]h!�4]�B�����Gmzɢ*uu��PM�:ׄ�s��!��^8/F	��W��2>���B=ӎ�C��KÌEOc��Nd�����������f;{#{'�H�l��Ge}3J*��;���US��?q'��>��<^x�C�|�-4�DRv-�KZ�K�CHT=�	�A��g��F�]� _TVU� /�	I�#P&�M0�E!��_�����{;ʙ,aD�1����C��0����l]�q��i��w�CVN일eHCLl��|�f�!%����M������.t��c[i0�g�s`�^����ϣw� �������k���y��{������v/W�w��ҭk�`�RX,�蘍9VOL�#�.	5��7���3m���a�����9�k>��˒�]���P���w��N�}4%�k��vԲ�^���x@�Qs�5g��x��Lx��v��pj&��1^o.猖Bߜ���,d����9�s��\���-��l�'	�U|��U���B��rT)C�		�}8��&������:��>� ��� �x���oA� �(����@��v�Lg[�G��d=�P�^��A~���%ȯ��G���VkOpt��/c�+�z���u6=����t�6��(*��%8
tr� �F4	�RE�	D�0�c��x���:�\�M�ic�
B=���zY�zY�8�/��E�g���	�N�X��4}�a� �W��X�J���甂x^�^�Eg��<� ��6JPL� �hϋ <���P���'@4@EA�ު4�7��U��gT s
@e9�m�} �V�mx|04Ia� 4:5R��&9L�˺!#J)�����fD*�(c&���Ϙl�kn�R7	��O�����Q*!��cu��h��&�O¨�Ftt����®@�w�/<���O��BJc
��
�B�>Չ�C�()&��V��I��G�$@
X#:�_A�n@Fh�9QLA�3H�� �R.����$�J"�J��ܐ��"Di�+�FR]
B��F �a���|\y��<7��G߾jD���Ӽ���[e,5��8�੃CA�s"�Ap��BBMN�ޏ�޺�����S]Ȯ6ƃ[v(���aW��
5p���K(p^4RKbQ^����D�D��"\�ژ�:®��b�8.Fj�:��pso5޻ԋ���A#�R��	��
�0��}���rDҶ�Ȱ_�>cc�&T���e�\�٭B$�a�|l��ץO���7�}@O�e( zu��;���6_zw��	�o�kQ���<{�W㙣�xn��L4�>;�[4 ��P�w�N>{ӱ�%�k��_g����7b�ת(d������s_I"�+3�V����$T�&�<'��Q(Hա�,�=�8sb/^|x_~�|��7��s��ҝ�x�:a��8N�n���z֕���]��h�+@]m.*ks��^���LD�����C�\3��;��5|O��?4��/��?������ ����)��X�����r�)X��
��#�#jY�{�+/��w�kv����}��yo�Á�n��wp���p�k��~	_����#�>��/�{�3�;1�h����Ü&-f�� YD%�W�����Y������o���_q�/����	����џ�,����xX?@Y���,'�S4=��\���`s:T���۞@?�]�O��s�X7��1�񷢞��gv�>�)���f��+�{�n
L	���{P�	 �K ���SƂ.�7bIO�FaEC4�[�ؑ���Ld4�{W~��G��_��	@|I�=�O�礦;~�?s�[�����W��{��7���&��C������� �yX՝�eiXN�\�+���.H�	�}B��\8�񘊷t�X�g�r�#�/�{㕬T�/K����F�����X�,YquXҨ��&.7V	���P��ViaE �$(ZD-	���.S��%|���U^ ���Y�x:�3"�)�`��M�<\�0�+}�3�ږ��s'w'AԾ2
ֹA
"%��q��K*�ݙ;��;�;��l�R�G�c��	+��Э�I ���0ϼW�Ք���,�JN5"��Qp+A�,v�ؑ�mF[l���&��)x��o�ϵX��7Y`��.� ��@8B�
�]9k���6�;���cK**'�Q|���Y�l�N�� ��9*LJ�,O��P�E��4�B���S��Q��Jdn3e�s*� *�8�����,�9	�2w�@{�q�0Ȳ�V��P�S�^�&���1�5� h5m���\�Ѝ���(�W��<�l������>��ZxG *.YE<�"�uY
��������oGO_R z�*��S��9r ��#����`BpT:�����3�KFPd,���٧2�8w	�>�S5a(*.DB\,��hC�k�5@����/�m��l���z#����=���"��G���[h\J¢#�����+ׯࣟ�e����R�Uv#��_�����_H�	���E(,i�!�ω>E���1�=|����w��cj�Ћw��/�yxna����F[,۾�-üe��{v�L,ݲ�6hjx�w����z��v��o��G��Rp)�9����P3-�r���]i�&d^4��9]��3M}��7�	���:�}��G��3Vc[*�3�g	%/:Z�b��x�f����R�[%|_T�D�J�� �֝�ƌ���P��(F	�c�/	���#�c�� ���7i��4�kRsG���֍����&�]�Ɓ��8x�W��9 Ɇ��	���4�T�CC�4ĸ@op��2@�|�����*�|B:H����1Q.��NE��q����>!z\&�sY$�!\�pBA/Hb���`�������G�D�sx��٤�,�B��H�4����`~~��2��( %h��Yr?�_ U�T�3L�u�W�ϧx<}�@�,�S���0r(%��A:/���(W�S<����PS 4q�,�^PM)Í�,Ӕ���9�RN�x>�������4*���t��	/S����O�0jȒ�CQH�
f�f������T�T�P�<� j��\��$����,5YQ
B5��͊�or �Mp�9Å�e@�?�kbQ:T� ��X3J{�Rö
�a,�@l)ϳ(� �(v�:��`�J�o:%nlI���E��2=� ��g4;�(	�@cJ�*󰾌�Y��pI�T�'��"(767X�ݐ�]������}8y���H14�p�sdBI �x�S^�r�`�
��冰�t��\���7����q��̭��4ٛ��}%s��!'���Xg�����*ODqj8ګ��X��Ԅ@yo���و�[��xWhO�;W���v�J��N#N6Fbo��3]Пl��8;京�~��(�݂��Ht���ێ�g �u"�v`ǲ��d1�+g!?�	��z�.�Q��]��F ������&uk	^:V�7�~z�*sr>�W�!��cu��J\g�~���ѾL&x�H�>�#U�h��AK�Z���I��L�B!+�oJ��5gD�)+�)�Ȋ	A���@�'<���1�����w܄p��\��1�1�ȋբ>7	e��(JGM�����0��E 73����ɋCYU����O�sd��&��|O�v�6�+S���S�x��7��W��w�}|�w?F��=ؘ�U�gW4
�%��V�̣��㱼7A��4��~o����?���������Ə��[��Ͽï�������"x��_�������� �޾���}��Ū�P,����V~^�Iym���\�~�_������).�� �޼�4R�O�`K��.� C�yB
D	e��38�Դ :%B��J����K��?�>��y��b�Ox9EO�fvROS�>/���I/��="��(����4�Ü�Z��O���|B��"�ru�����szc(��n�dyv�s��"n_���-�v�p(@P}�+R1q�,~��_�|�ÿ�����P٩��OI�}BO�甦;�����"@**��?���`��%d�T� ���IG:�7^��|��ª�,ߝ�e�E��"8
d.xB�]8�d�I���=Y�	����D��˹�b8��|�27�xA-��&,�3�����V#Vu�c]w����|�	�
B'��J+B�!Ԋ �@ �4�
`A�ȕy��a��I�h�yBg�:�{�!���dC{��ݩ�!c?	�6lW<����l�Ca��~�!����[_7����C�H���6��Vh��䂅Z[,��aa�ʹ ���*�m)��{�
E|��vg"����P8��6�6I��a���(l�܁�![��w=V9���f3��Y<��� @e���A���]<K�/VНA�� �� $tfMh�J6� t�� Z7	��
4�2�� *���b��XP��_�����d
&�U)����0:���N/�	�7:�@>B���A�^���&!�uW:�T$��?h�v4_�E˥>�W�I�٫����IɈMJ@x����^A�t�E@��ŵ߇='X��Sq��M��@��A��n��w"6�;]��죣-�SZ)�*ZU�g@$���0<~�o�E^q9�v��&=�3����G�5DPa��������*���7<��	W/�PI�֬[;[�MF$��"B���m� \�q��ַQPT�@��-�����)pp��Dz~�t��'"8<�𙍔�2�ա�k�/����^IH�������8|�".������|Oxc��#VZo¢�a��� ��f�r#�U(�_���-8���%�
��^�D��9>'��
By�k����
�^��ufy�Մ��K�*��!�T#���&�����:�㏵��@=�FJ�Н� 4m�@�e[L{�d���X��;ۂr���+e�	�G+���Z{�� �� ��%�>G }~
@w@�U�L�2��y�� �n���7c��&t�f�݇������������n@Mo2ⲽe	n��1� \:�htC\�'b$[��I%i��Q�h���o� �F�IP� ��E�(�r=tjY�R��@,
�� 3���e����=|�m��B�xS9N���l�����dY�S�T@4���sQP��fɺ?�I�s]`S�ԟ�<��F�'T�T�3��U��j���	�m��)��@Y
��B�H�sJ!z��@j�P?��4K���%�J9%�O	ՕP[��ǽ�a��N��u�JH�xEվ��}�&��tj]�@�P�֤t�%��� �#�E�Z� J�44WӐ�JY�ˍATJ�T�>M\7�Q�1f/��h���D�E#�* ��AXf��|�ŗ�d1&���"�>��(!�VJ+����1�2��U�<�C%0J��Y(�T	�\��@E�"�)}�ZL�%��	�ձ#<FE!��V�j�A����O��s8}�M=Y#(9��b{";�vʄ������#��H�i�E�"�J����;�^č�8x�Y��I��KF l�C�-7ֹ���f] �k,z�4�����~r�����+W�gk���X�La�Q�僋��6;�g�B�)Gj�0^艾TG��v�>b�[ z�LT��a�׼!����ZlY6���N�۲t6�}��s�d�n��h��	8ݖ����5����q}wA����k����f�rr@U���J�;�ȯ��?=����ho&��g�d6T��-�·x��,j'*uv(ہd��H��
�;����Έ�~��p݊0���zl��m#L^�b�����}�B8,������ݾn,�,D��&ćy"2�A^��wD��z�?� $&k�����L��梨4E������&oxg�#�� �����o����
��������擣ؖ���_W��aiO�
�0\J�ֲ7��ð�-��bϭ�8w�<>|�M|�[_�w>�6���?������{��/�����x���p���T���������� n5����,i7a~S4f$:b�����?��oq���0q�,���h���M��W���Cz��#	�N��Iϧ��ǠF�zBӃ��q���#�}Lӂ"���I	l�$d?.	y�!�Oh�� ؜�@���OH�R�PJ��ڔ��Y :��GY��5��O�G�b@汌���(�u>��i΄�>����/��7��<�C��?�񏏼�ӊ0����O�t���O6�?�P	�����78x�r[+Qd5�v#�H;��Ú�z�sV���c��,�P�'% �(�v$� ���㟆O���.#�.�'HR���Jݹ�O	ŝ�F�谈��.>��X�gM T���P���WM�m�t@痆â4���B�g��/�e�Ӗ�w4/V�~�H���TO�IpŌ�X����<��é9;٦}C��Ԏ}�gu\#Zf���&���7p����U�β��
@���]FY��@]2\�W!����($�U�oC��<h�~MZ�WV��`��	��mF;l��`C�6�؀�.+a�y��ًg���>���@E�.Ɉ>,Z �%VX�y9��m�m��e8Vz��
�-(!h�xϬ�EȤ @�֣�X��)�|RS *�)R��z��B��H��"��ВS��z0��oF��h�ۧ�����@  /���x?;�\�Q����[�*ޱ� PIR$P�拽�*�m�+殱�O�?�r�	�1����Ƙ@���g �I�(�n���>��9���q��;�}G�`h�QT4v#����<ڥ�3�#8*�vpmfB�d�5`�'$�����W�~�9��	
"𥢤�ɉ�ІE &2
����􇻝+���j�O8ں���9Y��Ķ�����FlB<2rhCEE����A8v���� ���������s�e]�������%!>��Qi��d�`�V����F�5�$K#N`��8t������b��i�z��x	a����VO'�ڹK6�]�PM$ :g�S�F��:T�D͉F%����# m�٧@s
>�4U�i(�]!��:�>k.6�o�F���@�:psNv��T����}�Ƞ�ԛ�xڛ飅�[�b�V���:�V�l@��*�,E���$��LTb�ȳ�#��??��wa�s�q¨d�~0�a���&o�NޠݼA��E�=���6b��6��|/-*�]�£ht�m@D�f��w"V�
c�+�Q��G�@�sA��ZJ#�;C�Mi�\��|L���H'�t���BX|��)�J��W
$4q]�S�p�_�^'aS�g�-o��m�v�T�,P���l�yFb��"	�5�	��]��H�OA�$�>�)�eR��}�����
`�T%�6d>J�7T�'��mJ�m�V��u�I���}B%�6P+��� ���4+@yD�(�J��)����)o�H�Kh� �����1�}j̨�M�#Qѓ�̺��7:=Qi�Ф�!25)V�Z�ЦG":S � �k�Q��C,�3�����X���Ό�6C��.�|y�67��QˋB$A4�@G�#*WMN²����x7�����	e�5q(��EnG�y���dZ2[�n@Z�	�� 	�&�^a�H5HȮ�i��&u����V��-#d���P]��Y n�v�6*�)�_=�W߹���Q�'��&;ؤ�#Nv�6�Wa�L�x��\��P��e�8qc��|ׯ��D2K#�fp���Mf0��F����/�-�7���5��*�ͷo��x��8�X�Esg�y�%2.h/	��=x�/��rq{4�[#q���9n��@g�
��@Kh5l���3z2#P����i5�-�� �-�܆�Kgb뒙p#���۠55y��ŉ�x\�I�ա,\��5������b�o��|�/FI$t�/���zcO).��4��H�@��e�HgˢPj�Gv�doAA����m(�pA%�纤t&a�:c�E��GoY
�k�q�� ��p�5\>�U��ͅ���`ez+r�E��M�"5e�g[Mu�h�jkr��\���
4������ehh(DE}��S�g$�Ȉ��*�y�^���~�&(~�_CݱAl���2V�W��=��=q����˃aߛ��ﾈo��O����ￄw��*�}���z'_��]7�����=��O��N���	�y������}�޹��s#-���̯�܊P8�ea��K8��}�|��޻�����sWq�[�w4��1O�;	=�i*WyB�C7-|�D��9	YS`����
��|��Й��z��z��8� g�v~��NS��Ѷ�E��'�>�h���@��1������%�3�b`�oĲv�2ԓ���t�6�������w
>�>F� ���gU����r�Ok�������?�G�N���u�i�D��A����l�]��{�rO��g*�|R�	j����8�U�,W8��r�!3t.�2t�@����"�B-�L��+��].ḄЅM2?��뢰���y�xA��� ��@-��[���y�EQ��BU�ܕ5�X^� T�O�¼dXD�$�`n���z�7�	��t��MF85�RC ��)/�%:�:;�;�^�������S�����]y@e���(;,��7?d۴ *y@�[h���Q~��p5��cEЍ�"�� ��HxBr�`�ꂭq��l��:�6�ڈ5���`��# ����)^��	�s'K�* ]�@%� ���	�pl[23�C�
@K	��t�q ��,�h ��'��5���@�8�N�ފ�Wy=�,R��C
>e�xA����#xa�˒�`y�MA�,7^�P^O�O���B�xƦ��K�	���yBco>���@@�bDC[#!��RNL)�������b~��zTֵ����"���{p/:��U\SZ!bӋ�^X���}�' � ī����[��;c���8�:��3i��3P^Q���d�&m4��a�s�3�Ӎ���C��z�-|<��Pׄ����������RS�����38"z�����o���:����������-lAPx*� ������2D�3	�Y����R�<�iy(�iA��#?r�����ӗ��0����N߹����G ��v�mY��k��j�9�̥3��oR�d�x$|�{�Zo��Zn���[�2������h(�eh��z���D5��4c��1rw/�&�	��h:ݫƀ
��we"�/[�U!��c@B+��;�t��}�	��X�e�����=X�r���Gq��y��]���8�<��G^ه#/�c�n��(�o�c�7��{C8��a���?�{	����P���l	1�Npۄ��M���
���蝈������p�#�鴄P�iipFh�"�D]��HBh�	�1��G�tR�.�dY���,��Lh��PY�:�Η�@�x>%�6T��u������[�'4D����iQ���G���l���*�V TBtdN�I0�N�yI�:��z+u���vp�����x�Sc?pV�g�����Po~G�)�@%�o�+��	��ƄN��WT�{�>�A�,��))'%c@�����T ��q���vY��) ����FE�8Q�&CK �1���ph\�#<5!�2Gi ���o�o��W�v���6Qh2!U�!\j34lC��PPG �-4!��x���c�e�W�����C ��+ ��t��hBh$!4$;��x'��=�n&7x�{�3�ׂ���(��$"�3����u(��C*��D��4	��ݤt���H$U���"�@cX[#�+!�s	�%�Hk�@pa$v��2`��/�"$�¹s��b��!��A u�p�u*!4��������u�+�3���@��CϞb\e�r�R7��c�๸�ma�nI^��0�H� L�BV�-��8y�	_{�^�3�̸ �X0�΀��*��c�F�3'�psw.n�X�7�����/rG_�3�S�P��A��r-��+����j�g��J,��o�Nx;o�	�]�4�W�D��4%a _��5F�h�ù�$\����l� ���[L�-�+'j	��xM%!����I����b\�5;ڞ��=�4��pwu��@[2��bP���i[��)>���ZT�٨�Amj�rLh/H@_y*���ڞF<s������x�h�=օ{G�[����`-�����7���˧p|�NŹ�{���9ܽy�n����ś���s�^���_Ńp��n􍶢�1�"���(B� �1�~�~����k��!�����p�.��r�gN:$�Ldh+��<�tz����_���#|�'��/>��3�0�gó��X�⁵9~�R
�b#�v�#����/��_���������q�_TSX����S�������o����	�|�5\xp���.�t^����(�21�	`S��y�y}f��`�RIy���09	c������'������>)�^J�$�$�}R:VՎ�-��Ҍ>¤7@�2bΈ	O�3Y�����cMWg�쁘OI��i����%�̚M��[�f 5a>e�K��F��Ǆ�=�+�_U"�5�8v�<~���H�3����*����E��̷�W��=	��s�d�cz���?���p��YBh=�&FQ}qR��w5���c�hV@W��'\�<&3���SM�"�p	�\�r�H*V��a��s,C���|�\�fw�Z_ Ӿp�����e4g��0@�j�xA���Q����%�tL�щϽ�P�&
V|�,+"0�<�	���OP+B��TƂ�����,_Xf��2�(�t/�0Yc��닃�ٝ߾��WIB��>�6# ~��=5�g޹C ���'�)����?�N�"lZFX���Rˈ�*	�f�s�rB�Fy�O �4�#�7���~o'J�K�f ���𬖤y�t�wdB���c�Vl�\�%;a��Y��T�`!tJ���P�Ϲ�s1��9g�̵�:J�G!�� �� �h�B,ݸ�=��3����H�!g�F6�� �n�eށr��( � ���t�6Y��S!�f��y��9��	���?V� 4�ea���1�	��[�|*	`H^lQO	���v+@�v�Ɉj��t Zw� B�h���/��q��=y��m��K`ʈ���p��*�	ٕ��2��3��U
S"�|�Gϩ���ڏ��]�i�GqM�r*����[ڌ枽Ȗ��I��e�=0
�dL��������}�#�0&Pu:��a�3"<4�^j�X���p�����*������T�>~�ȶ��ŗPTR���x��N&�ư�֎V;~]��-�j|gRj9L��HΨ%h7��\����%�\��UnMS��;�[�kZހʖn��~_��w�����]���s�}�4�
���m^�
@�o]�EP���0��)�^��hS5�C!��XƟ?�=�L��� n��~<���IUʔ+�,�Bt��r�U^W�����iX�'*��������O�z@O�[��8hBo6��x�Mfv�1�����|�2Tೊ����@��25���Bp/�v7�p��?��_��L��q����N���`y�Ӹ��.>��~g�ۃ}���:����$���&�mDP�&��mEd�v���|��F9@O�=-�MC�ҰԲN���=B�����H�j��3��CE���p�hڱt ��B��tU�)�?E
@8P�N���P���e��Gp 麟�F8Q�?٦��<_�
lz:]�N����+j_���N�cRP~��t
D��S�R�p[���������ם0��sP����V%�����O�x@� �O�)��T^�O ��Gy;#c�!�2�3<������I�|>!�)�T�9Y'�S��@3�<^t��)u�)���o')S��H�H*��J�?�Ɨ���O�|��$��(%D�B�~�m
T�c	Ւ� � O�����O��=�w�Gr0S��hh��ل�,B_f$"�#���|��������+��)6�0���=��4���c�ˇ��@-j��Q؝��ZbJ4бS�OJWh.��)�
ϕ��H�I�m�1eQЗF�D�y<��i���7����[*�9������c��J5���?�� ���g�=��;`+!tK�6���:n'�|F�<�1��������a�8�αR�8������ؔ���}^8\�����#�&�MI84Z�7L`oO)��V`5�sǺ�q_��8/�'Ľz��v��l���±���YhO�Gs�#J��"�n��8�Eh��B;�Y�\C��X:W �ρ�fl\6=�U3��Ɂ(�b?A~���3��җ�k�Y�>������;��9�糇+pon�#�B��"����H[F*�0RkP�|��ڑ����UbpE��Fĸ�A�I���M0zn��{2"<P�{���@SV�7g��H9!���P�s)�E��iv�G;s��9����J��޸����x��8zpm�%h�+@ME&:ZJqho/����pv�����p��	v���:܀̆,D�NLm�C��>�����ڏ���M���eT�}a460%	тN�$|Z�0�9
�K���\���/���#|�����w�v���V&{`Q��b~�/��`v�7��ñ&�Z�ui� ;@Ŀ�x/~�M|�O���?� ��J,L��U�7����ÿ�_�շ��{/����q��%\z��B[/�ok:�Kx �BA�d(.Am�$t>)�p�L��{?C*��sH<��OJ'�������%�@y�
>��fROK��4���13�O@g=���K tv?!��j�0��f����"���<�P�c�>�)-�ú�D��*Axg�k2p��Y����nŧ�w�_�,������t~����\ :������������ӯq���vգxw*.�B�^�����B�ߕ�ec�*�v�h*��TBp� � ��,�Е�X! �+S��S@�x(YM�"Y��t�T���Y�p���3N���x��m�XB-&�.h4`~-�S T�j-,+#aA� �Γ��qs0/?@�E�,��2G�%o�Os�L���S�OTiU2"�V���	W^L��H�����}ϼu����>��nX��W�%���N\@�\�݉��S�sC�F�E"�����D$��d:�!�tb�S��4�C��p8��.��i�؞l��6E�����X�s�y�9����I ��U����9��f �0���N��'t��� �څ�����V���<��G��Je��<�)#�� TBp���T<�S�QY�DC�����P���{�s����v�O����T���K��V��Tpo 	 �W�H@%�gh��N5�d���>�SK�{�ź��z��5�:9�%H��G\Z�	��M!�e���g�c
>[:F��/��w�B��QԈ��T����Q�9�OS	��8u�6~�Q z�������ĴT�f�!*Z��� �ш��"���ށp���N'�P'/�y FkDCu#NB_x����!++q	�p�����<�;��ΜAK[�J���Y����}�U�hhۃ��NhY��x��|�g���;d�W#1���،T4w���[���[8|�FUYp��E,�C�>�Xk�+����uKU� �e3H����M��F�+ *c@��^�\�~n��>+x-��P�@��=SI�j�֡�pXE����A�ك�#-�;�Eu*hޮ
$��) M-Tsي�_<���k�֝�}#	�ζ* -�* *Yp��u�r7�� =H����&�OԠ�P9z�A.��;v���]y[<��4����)�	�>�I" F[#"چ��<�J��:g��0ܠ��Mp��F�HJ�ڌֻA�B�$�j	��
@���!���Cm�d� T��x�y�y�PB�Ը�� T2�J�[�xH��`)��!vp��
��*W%*b[�Bp�KJHu��� k���;U8��x)4�� �'қ��T
hJ(����OK���<|$<X�I�˲7���)�9��V��"_�'ɉ���
d�!T<���[��9A>U(���d����H�%�6�hN:��� �qM��XJ�t *�S�>��s�@T�g�1l�(`*mų��`�(Ż�8��=�<@M� ���T�����@���+�O�<�n�ߍ@#r1z�)����t����ϋ�gB�5���Rh2"�)�0�<	��9�IFs"�z��������b]����4�e����T���ezs�ؑJ�[Sy4j�H��Qa��1��
@�X� �QhL�����P�M�Y�� l78�wCZc2_���(@)"*��E�l��=�[����%��Xn4�`��6ڍ�dy�oO�_���ό���F��0	Iv�c";�� l�
Ŷ��@���4@j;S�Օ�q��3���a���X�d6χ��REZ(�e�͋}��b�h�¡Jf;�-qb�Qg�C��fw,B04�v�xݚ������z���X#�m6/��MP~��y5Jx-;2�1R�U�8�d�ŮdBh�����H��!��)Ľ}Ÿ����ށr�"����H&�}v�0L�ios>�vg��Ʈ�d�$�#l�x���(�5лmD��rج@��z�9"��Y��Mّ8Ҟ����<��[�E�Ɨ�Ł<��}p�3����Q����䋴n���~�5=4���x�P[��c��qxO������g�w��J@$ӱd5f�X���2#ܳyO�q��	��?~�������w�ǉ� ��ּg7VFcY�$pR�ȢU��E�XS��gO����-|�����;��?\�54���cI}$�D��#�<�F�V��V�AX���&n��k�x�����w�A�X-6f�`KI�J>4�8��=�z�
��9�s�^��7���7�|v���X_�#̘0��# *�)�>� ��O�x+��9��|ғ�������Z?�ޞ� ܴ �s�4'��׌^µ f?�G�
� ���z��8����94[�|�fr?�=�F�ٔ?���o�5��i��3K�㱦+.C���BX5��F�����S<������������Ѵ�ȿ�@'�O�3�]�%����?�.޺� �ab�7�@w�.{ʱeWVg`ٮt,OW *^��	@�r� � �� *�R?���Q��s{	�]1�j�eT��$�UF��x,�5-�S��9�ј[����g���)Z敇c.tA5a�4s
	���*
VS�Xd�a>e��J>X��E�xڰ34��0�E%"�\��(������b�1vz_�;��/<�4�2Y�A���j����e:',��Fm�,�ے��4,���J3�&��t+����\%�w��H���ܢ�gE\
}`�펝�؞�m1�p���j�����i�Z4{@-��t�֕�񱅋��	m��B���נ�P���Hn�d�%HNy:����� *��R�1l>���1@s&T�c�q���	WM���]iE��f���w�
p��S�D����h��>�\�~W��}�9M mN�6{<;Y���W/�oh�"��GR	�%�O+$����3�ch�0[1<~�,�I���jUwa`�I�8�Ρ#(k�-L ��H�}��w������;�w��kk������d�''@��Fc}=�_����f�x�t����\l��Kus�@�o��à	� ,0:��)i��bj4����\�t���/��o"JgͶh�څ�~��ص��S*PXэ�G!�qI�HN/Clb�ʂ���Wpm�t�ס�{-}��؅�GO�ԍ[9v������N�w܁U;6`��e�\6��K�G ��D�/�_�Ğ�`�+��qg�����=������:U�ʉZ��߫ƀ���V�Ke��$D�M�}�Л�4�O�j�#U(!/J�ڳ-h8߆�K�(?Z�⃥���	B��R�КZ�򃐘�C�3��f�EH!L�!T��!��	Z������^��kK	H	@[�|�6~�	P��iv��({F�4!�K�$F�^�L�&|����	�5+0����!���Oɲ�g)�~!;`��O�OQ�v+:�
hʸ�ǥ�{
 *�*!�
JY'p) *���1��
:�n�=���g�-<w�R`T�tʼ����
|JX�WT���;*�p	Pr;����[z+u� :��S :��|<�<ԇ�RJv\�Ox?� ���ƀ>�)�TM�O��@�d�d]%J
S�ǐmr"��B �7������n�q��ol ��~�&(��/�̀�`����B�T���Zh��c�:���N�$�r5J���WSO�#�$"��e�	���E�P��9a�!�E��Z�c�`{Ay����{;�D/x��tK��	^�n�" ��@W�AzS2r;2�ْ��$d��#�9����j=��5�* _�S * Wm��"FyA�ez��� �(;��ء�'Ěp�� ._���b��aH��gx���f�Ɩ؝�P{�6�'4��I�p��m�����<��ء2�#(�NI��
���X>��i`@����{���w��D+��8���p�\3�Ẁ�����ު�Nt���K����Gh��+�C_�=�㷣�\���	�-V�ɶ���������0v;�b4�}+¼i�����E��Cƅ�X��`Bl�z���$���8��]2/h*��g��h6���W ��@��ޡ��"\+��,nM����-�8Ԟ�#�y8ܙ�ڔ�o[ �5s�q\�HBg0KI4���A,��d�t��yojM���\��3�pm�� ���=��$UP���
�z�,~�����70�ߌֺ��U���>�BqV,��v�u�rl"�Z�n�;���X;��S��P��r���=��Ͽ�����毿�w~���%5�J5*W�9�&2�Lƀ.ohI0V����!�����_��WQw��	�kyܲ�8��#�PsM�7O�:	KیX��"=v];�W��&�������4�5?6�]��
���{�h�5�yb�޼�׾�|�%�ѐ$����&�|~ ��9�S��i�7N�	��,) 0�<���A��z� �d��ha�)�G�YRӴ�2:%�vpz��t.��#�v���OH����C�Ԥ$����(��X̗�[��A����D���#|�Q��������|BBd���9"�#��|S�y4��t *�:@���g�q[� ����L ����]@Yo#�N�������'�hl�ؓ��3T�[��O �� �L ���b����Qs�"ɒ��0*�)ɋ@-��Ԣ��%s�.��^�X,'���N���V>ۍ:̫�b�@'Ԣ�e���s�B���糜]��Y�����y���?X
�R��|),����tw,Lv�U��gzaKI�P�#֛�actá�{�o����Ğӣ0�=����PP��e	��ń������t/���(��7�6����l5����.T#yO:����XDv�P�� ����j���X{���\�Z�̅3'Cp��tնUpt�7m'��0��������]��&��+W��#�Z��<���S�@�P3�~���2�J��b�-A�Z�2�L�"0�H	��\jQ����h
@�ڭ�|��� �|��@[����J?�I]9��Kf#� w��G @LBb�h�:��QP�D��ɳ7�շeU<��1T�v#-���}(��!��ƾ��j��`*I�2�k�^X��GN������;�1�g/r��������l��H�v�
~���`����p�F����m=8v�8�َ&Xww��� �'aA�HKNE^N.�z=���PH ����w>��~���H5��eN~�qE��|1b�aJ*�ޔ��_IH�6]*Y%V�_D�2Q�ԁ=gp�γ8x�����h�)/>:~F�68Yc��� j�h6f-���� t��D��n�]���0��~�+ Z{���@k�כ���l��30rw�Nw��Mt�d=2���Н���L���h�L���	��x-O�B�xA�.v�ǀN�In���B�ف��
�@(�@�ۨHQ!��a�̈���rP������r�p_���K��SBVR���c5����f�U�Dm�����6��`�;)'��p�O�J�۔<����w��,�Y+��ܡ�{l��?�d.�`��$��t *c==��9����x3ElC<��ޓu��1��A;�	��2�S���K�<�ϧ�s��@�xCel���P­�(�M`U�T����, ��c!���S<�f+S�HحH�TƂN��~"wr��9���ǂ
�
��k$Y�,���N�*�B��_�ק$o�2���e��
�}<�Д��U�D�$����R_���}|L,	��^F�xM�x�&�/�pJ�K��T��d[`j(�>O�88������xg�sL�gF<Xz�t'��gj��E!98.Dyc}�����W�<��{f<����'��H�GJ ܒ|��ePv�nI^p�s���Ye��f*�iO�ZSQM�q_-jwU��7���H�7!�R�Xv�	�1H�5!�>�U&h��.�BZG��a���xW$����Q<��!\9׍��<ĥx�C��cm�5� *��Nx����a��?B�O�+t44�Fsq��CvD��!�(��ߙ �H�-����H	�����o7^{p� :��(l^2[W>�-�!�����k܇/�c5:��z�#��[Q�U48�=�#|��@m��:�U�7s	��;�a��i�~4&V-P j�l<6́�c-*b\Еᇱ�P��©&���s�f�ԗ��C��9��[�
psW!n�.V�ym�WǋU�S��mI��c�<C�1�ݔ����}�sBlWB�N��w���ylA8��يL���0Vc���X��J�u~���,���ĩ�4��6T���h4h�R���$������-��ESy6�p�]'�5pq�7��p���[�=�"��W��S��9ފ��%�6h>1���E|�;_ķ~�}|��?A���� �)���V��N�GP��,[�_��4���9�o��{��?~����;�4z��0+����;�ר�>�K8��])*iʊJ-\�M�5�W��.^��{����:܎5�!XS�W^��aXY��u�c����+x�G_�ï�����"d�K+#?�+�>1��iT�( �����I��,	�>�/�I)`$,>)�O�S0g:��#�4���M�=�c>��f�s�>�b?��)�Ü�X%9n���투>���p�� �?\���B$����k���#��)���|���b�ϩ����O�ԟ����L�"���,u�O5,�3ç�������?����(jAӍÈ;�͡2�ڗM��2B�@e*��@	�� P�ePY�}S�T�R��������b)��wi'��L��s;�>
s	�uQ���y��S�9�%��S��E��s|0+��������WS�,����lh���ai�'Vdyaq��
�]��
���wK���p��!������u���YZ5����t9���uf �r���&�*�}z�V�L�Rq��w��B-Rv�#� C ��ApC$|+��^��\O�L#��s�r�ЙP�WQ���<wŖp	�����H��Y�Bp�N�(ϐУ�Zɂ+�(e�D�
Ý@��)!��%z>E�%|N�-?[��S�p� tj*��+mO���ǀJ�[IN$ɇ��?kІK�h�އ�[Ó ڍ��"8Dz���s�����n����(��ENI%*�:Q�1��^T�w�����}(�hEy5ᤦ}����UT��">�2�6�p�����z4t#!��e���#���ߏ��b�5M�H�JG�N�A�_>w��E�s��fk����O��G�������p|�q�ں����BCg4!-%��H8;;������_㗿�%���O��B�K@DT2�"�2ߩ����`M*�2�]k��Po�h�i��]���n�֡��	%�m�ۇ�箠kp*�;0t��O�DN]��я T<��&Cp-���\�4��P�_�E��n�^���s�6^�W!�2��)�N%!�=ݨBp@Ou��8����l@4�3�]�H�S jÕdDU*W�~V�lD�fTL�<��E��R*7+�9	n�O�A^�/2�����	1E1��39S.0q���&|;��6��o!s�;-�zץXK�rZ��K��a)��-�❋��Z�s�Xa���k�a��Rlr\��p��瀭p�'�p�� G��nka�;]V��m��6<���f�zm��7�p��G(%\�
�	|���V�l	y~�;�F��X۔\؆ȃ0+��F�u�vW�������=�Z�j���<X'�e¬+!V�\	�nӀ�;a�=�4 =C�d�-�VI���;��I�����.�⺇���DX�p	�u��ղ@�O8�)_���JB"������*I�<}��-���4���'���yxf�e_�>�Y_���S�~:/��Mo.{�NJ_©Z�1�� ,�j�������8.�<��J^1�NO�3�G��t�񄳁P�s�}�����:'�9�6�'\L�p2z��u�۰����k=��n�Rj��,�^+�����y�-�؀%���n%�X/��+��~ֲ~k�N��]`k���hXK���F��Xogr�Nv�6vv"�#<�+�g����I�tBvf��R�Pf@Zs�{��e�/A�@.2%L�BO 5"�p�\�N��� (a%�=�|N���	��-���x�� ����=eH�"Gm�]�v&8aG�#6�.ƖF�;�@DT�C/�� =#��}������()'���k2_ ��:ؕ���sv�ϳ7�;Sp�t+^����T#�s6/��m+g�i�B��mP��K����>�v�g�Ⱛ�m�֨5lFy�6�F� �y5W�D8�5��W�rދ���Y�5P/���
�wY� ����V®_ȡ�K�a�&����q�\�u18���2-K'�'W��q}87	�
B�pm4���qcO�
Ž2V�cđ�ht�Z���[�GE����o��M���9o@��zxۭ���28�F��&/4g�b���&k����8 ��3� ����P��ǒ$$G�����p$�t�6�#.�~[�u%<�7��i3�=����G:Ë��c�7�y=�ZS�N���ދ�����_}_��x�o���AѮflL���0,�A* 9�]�����5i17�ۋ�8��U|�������Ͽ� ԺR���%缁8��d=�Ǭ�$����Z�k�1�������G_��o���}X��%4z�x�ݡWc��HcvU����o���=� T;^�Ul�R�� ��xC	��'���C�d,�fR%c�ӄQ�+�Z�n:�~�G*	ГIJ���r
պ(��� ��94������� *��)��)+zZ�u�IژC|RsEC�����>�Y��YÄ��4[�'���'���o�O�]Y���ϥ��>�	�p%Bk�Qw���;<��������_�L������ɂ>�o
.?����>Ej%g��I ��_�����I���{�T(n���>�	�'�w�t�h*%c�@����|����`.%�
�J)й��)��S�K��Mp�1�����?AE2Xu�yn��- J�j��E�s��|�:�X�j0�&s��a�]N -��B�$�΢$wn�?�	�9A� TA(5�}�"��R./�h��o����R��D��caFN���[���[�p��I�
b��mI�X�~l�� �wVI�jl�Dk��w��>���>(D��oL�C��>�� Z��}YH ܛ��1!�1~U!�*�k>���	�p�q�*ڐO����h&�) %P>U�!PK�vK �L@$��)�TӰ,�R j��
K7/�S�+4HhHA4"�L(��w`v]���e��affffffff�F�H3#f&�ٲ��۱;q��$M��i�����_gF��q����������덇��{���������u|�G�!c��z��f��\L��~@�\�x�
@�z�t�P���:Qu���Qs��s�����#[0v{�o���(��}~��(�9|m
���T��ȼ0����K���Q"ׄr��I_���Gwb��=��C�Q3ߎ����X���xl�3����Csw:�&�>��M��m�}S�`�&�0<9���a�oڋ�'�ar�A�_��^P�ܲf��W AЗ]߰U����O��ǟ�c'�ST���vܺs�fgh�L�ܔ����DD#!"O�y�����w�������������d�t�����(-)E\|B�C�;Ћ�7�c�νHN���$�"!�X]�����	QrV-���u���7!(41	y����ȆyU�[GH�Դ!%���%�-�EiC��z��z
E�-�H�[T0�
3T�\��Vc��J�3[���T�^ن�+�������	�z�(�o��s}��}@/�ߍB(�����0z���d/:�������mXv��(w��92N��&�S��ey�xk�v7sm�~��}���q7:N��t�@'A�~��;�! =څ��}X�P�����8��� ���P^��� ��]��|&����,d�{"%��.�!�X��
0����!t|��kġ1t�8�4����r|��>ֻ�AߍX�4���m
W+x���Te��P�`+��.ħ��	�3���3ҁ�sV��������Z��aX�+�c]U�i�Ԩ��qL,���L�'�j��G��wC`�9�e<���N�K�ӏ�(�
8�K@�;�c<K����5}Ud<0�	N�SCY_�8O/��$D��ȋ��F���Ԇ��j^X�?�*��D&��		B�aq��@F�2L Hdy �D�."2����u?[���S�.&0�ϑ���E)	]��!H���BBTGC�|�t:�鵖-�D`^���S���8�x1ޚ�z��b�QM�m��� �������
_<�g��e�C�a��V{a=�Sw�� ����i+~�����O�m�l�>�T�%��cŁǌS�?\x�2�X��Px�n�l@a��S�"=���f��s-h�֌�ը(BQG6
����Td�&�z�
�U	�7��8��	����x�c�ss;��� ����𕎈
}�^H�P�R�2b��c¸<�2�D��3x��x��V�K3�$��ç1.,L��g"�'�����A�t�����۱gs-"�}=l���b<�����p�X�/�㩣8Â���P���;�-��h��V�m�X�U��b/sԅ����p��3ج_F��!5�nZIO�+�l����(�w�IxMVD`�.�Rp�/W��qm��'�puS��T���jܘ��M�H0����i.O����\��<2Z���d��Gb�,
-��bx��Z��@k��9"!���&#�#<�d��8W�d�q1�m��ޮ<����ә���TۭLg6&�30X����H�Ez %�i�~H	�A��WN��5���������0���ǂUI�*�a�ϫ���4h���(�;o�O~�c|�G_ë��]��#m��0lO��p:�Nf`�X�Me���tm(���������k?�:^��Wоu	�"M�`�B��,��y�'�u3|nb�t�nå�z�^�����?~o|�}=4w�x +��a�|1���cو�Ձo�������w���c'�:��4UK���YA�, q|-#�V.̓��R+�_�fbk��B��73���/d+��R��Ժ
�K�������0�|���/��9r��sY1�p[ܟ���l�"������ϱr��sYŬ&2�0����f�xZ���+��l),���ES���ǝ7���g�m�k��7�_8*r��@����§��OV����a��0�Az��G0:�	�E������FX�#$��KL�� $��A3��T!��"����v�&���ZRi�+׌��6���m\�=Ց��h�x\'�sOd���V������{8+���7+���Õ=�g7�E�v�cU{V�+[��� ]�����6k�M�wMCp����j�O�U�<�js\��uŁX����p��§,mSu8~� �z�I\z�:����SOdF�� &�D('ҽ�������\V ٜ���d���d��g&��},8��h�wU!��+cS�hL�zb�&������oeL�,�����[���k���T��w#��������Ӗ�R>F{=t�u�mXV묁��Cy^΋Flu*bҐ��{��tB��^�m�zP���h�T��5��k�&ݪM/�r3��P��8�0%4��R��0��Dh;Tl���A2���oOc��$o����u���0�^Bt�0t���Df�C��>3��3��{h�7��{n��N��<$�aٌ-�������qI����B���1�4��)�etͽ�����"l�X!J'�I�mڍ��;Q�>�6��|���*">K���S���t�d�#.9���8�O��g��[��ƛ�DZN�:�q��a����� ���!$[��Q�����r<J����kx����ѧ_Ǔ�=���,�f�app�\�������#lp��-��h=|�bc�OP���!5��	���/@f^jGQP��t`rz76nއ��V�fV %�\5ōK*Du]/Q�YuP�W҈����
��}����KO�sd��<`�j3h���uˠm��]�sk�\�����{�8�9���[�c}7�5�^Y���bM����w.��4��#�:7�������v���ư���vk�hϑ)"��ݞ~�m�T�a��[#U�|G=j�6s�nG�q��G:�r����yj���CQ�v�KEjD�OaYcY�L!Z�㋪�PT��SʂW	v2,氈���Gv�7�Rܑ@��JAh����xz@W �B�6�i{�����Z3�^&p��O��i�`k��,ԹX��pda���TM{���D#!�Fd2ğ4�]l>+�lU������t�����K����d(�P�|?�U����Td�":�Y�Y�+Ð/�N�P~�0��%@���rg<J��
&���G����~�Wy���
d5 %0CM�ɌL#>��E����$I���T ]D�B4�\ %�ey��NJ�dF0�9O��PΗ�p��eYR�B�
F9��Kϴy���)�K��"�I����p��P�S:�H����xeRI^p!:��}��g�S �,�D�+q����a�X�K\�+�	M�� #<h�eYl�ՁfX�o_3�������ħ��%���ۧ��ްN��B,S<`�����3&��0Is�i���=a���yܘ&��8�	���0Op�A��"���܁4�4�aS��*P�_���|2�9���E\M"�����Pڑ��f���G��u����#:�	���+�O�?�J�Qw�;�¾�X�q�_�R	Q�#�g�ܝ�vnm-�K�C@�/\���ؔ� �՚���,T��czN����ga�t5�ݴ�j�vƄ��j$;�)/ۇ�ps+.m�ı�T�j	�X��jCd�)��X �b-��!�A���$B��o��X�^g\�� !��.�07X�Up�_	kd��Q�ⅾ� La�&
��г�9�0T�scE���W6U�!z�'�s������i%@[���v<Ƃ���8�BΑ��vd`�*�y�H2G��6�͑$M��8�Dj��"�Q�j��f�{��\����t�6�bkC�b��%�-)�n��6���8<�c����p?��������Z������}�"�9o������Kq(��BaR��h���`e�/�yx�!������'��o����
v�â:JTg(k&�@�n��bTk�e�Ӧ6�W��ﾏ��gx�����-��yk,���"�O��dc!��V���T������sK�oǋ��*>��o�O�������ʆ�(QF譟/Q����KF�l��?|�~�"�8��-�0�[����/��������*>Ͻ��X
�R#(YĤ�'����'Q�hUm����@Wn+�B�§da���|@���ĦܷR����sA��0�-�+!釆�?Ҋу���K~��+�&�IϷ����X����>%������>ǟ��* ��������y�h?���Ó��=M0�S��5Dh%���fJa@��2�3R�)=�rzNO�y"Uz�U)_�Ȩ\5���z��kƫ=á\�=��z�]3�c�Q�k�	�U� �O� TB|.'>�w�aEG��� t��ˬm�)Z����.R!tuU(VV�b9����\K|j�:�n�e!�)�iQL���Y�������y<�γ8����5¿,	�%Q
�F��g�t�[�@�ZR@3GKP����'0��~�]EݱV��F>���M�HOG�p
b���[���`��Ç�y��	�u���@u�CW_���Z"v����)�[4d"�&	�<��@ڴ�n��B'-
��^���<�-W�Ж��hf�"�ؔ4H�'*�e� �l��g��.4�$@��S��؀���8.+��0zec׶`��F�^��y��C���ﻰ���s�a�����a�A�'��{�!�(#3��0���^4twcp�fl�݅��QT6�sw�����b`b���;�eu݈O/QI�d9&)�1IH�)Br�یl�s ?��_��÷��NT54���Օ��(G}U%��0�݃����Ԅ!"���������_�?�>x�C;|�y�cj�ϒ�rddg���=���?� �q�.��� %�y�̮At\>�K�RNL�;�@U�ʫ	��f��#1�1	��j�T�܊~�����Fm[/��6�G��ɓH�*����q������+��kк�	'�?� ���v~�,v>�l�w*��ؒ �f�K� �<9����=1� ����>$�� �e� �wt�h�9��(�R����hZ�q?<֍��
�]��|L��^�V�P�S�X�\���`4��V���L/"4��D(��rZ��\�,2X�NJtEL���ai즫irK�j�Zħ��!�{`���ԁ�~�-$ޝ@s���\�-��gN|�)|:�^�
�����k����7Lj?	L�e!j���)	 �U5h�pP���,@*�r�j7.]�\z��)L��}	^A�/_�'�Q�w��#߻��9�m�ʂ�=����\'�[",\{�:Í�t�G5��d|"Y�pU���Q�Ԇ��x�E�`t�6T�)Mg�|jzoT��bG�Ԁ�l��jC	R��`���ʸ��D`*� 4AN�s�B�$�q��T>oZ�B ��̒��,�Sn���:�k=C���·G������F I�XbS��$(#@Ҽa���PK�	0�� S�4�� c<l�e��`Y�	��b��)��o�z�r�%@94��e�+��:v�~�p�sB�,��s1e��a�����$��<�L�=`�eF�.0Iq�a�3t�m�e�Hs�X�*��in*E<|�Zӑד���T�V�iS#R�ӈ� ���f��/�������mظ�
��ܷӭ�/5��'�Fx�����<�L`e0b��t�tbS���M��\>=���4$�{ ��۹,�pmM�K}��Qؗ��'���;�߼�3�{�m������p�XC�٣!';G�peW�l,¡�$lo�0�ܑl��84�8���
)6Z�7Y��u(�Ey�������N|^+�e򲀏�),�V�Zol�V��t-�\�P�c����,/l,	����H���L�KSeDh.�	�k�j5 �ۆ[�[�0�Rz{o��.���Z/�\w&����[�fn��d��<�e)L�ʓ<QE|�mف�+�Hi$�K�0Y�����S܎�����@M2�3C��������p�9��^.�%:}�� � ��;�y�'��}ކ�;���A�1�	X]���g/��>��{��ￎ7�.F��Um;�5����,���b�D���`�(Q�;�vӵ��o����7x�ӷ�sh�c��c`5��r��,�pZ[���6�������>����^�W��!���k�;�E�zL�!,�:"f5���'	�;�p������3x������sH��B���/�^�y��?��p	�-6M�7+@i�zw�4S������$K6��Ȳ��?P����KD՘ޗ�����KU�A��x�5��*�b���;��%#��ڳ�a&���c��[Ճ��2���w�[
����߿i�, ���i��!�4}��70�w+�/@���M���:�ή*���D�Ԅ�n�[��D�������	<w��yj>�e�,�a��uY/�&�R{:S��Ҵ�����uo_��t@S��]ї�hO���JjA���Xב����8�o����(�&@WU�`%��+��pPm�S�:���ny(JC`V�� D4�b��&���x�/���(�APE*ܫ`U� f���K4�1I��ȝ�@�l�����nt]"��Q���;+���(�pS&3?��jA�!-�����4�JP��V{5Ay?4���淚�?�Y~e��ka��6lXF�AB}�h����0l{:�J46�kW�l:̨ZOM�R+� J��葁/ ��a�Z�|��|L�fTjG�q������)@�O��ⰂG��I��� W@����/ƾ��c�#;T'C�4��Q%T8�Y��,�LޚUHi̓��)JR�e�vه����ܶ�v`��c��٥�Z�:���m�<�ӻUM�Զ�/oA`d:��s�R��4~��%H�*DHd<��1�qF5��߳-]]�&f{Q^U���*��ee�4>��gϢ����	�z�������������෿�^~�e�$�������ThDT4
��q��%|��'^S5��a��ɭAzf%R���Zd�K/�ժ�m,!*�R��
��x�� 2&���U�D2�/jDO�&LL�D�tHt��^����Yĕ�	h���T_P�eз���!�}�6���?���]Ŏ�a�a~߷6�;�w�@��� �f�r�f��!l��{�>�.�
���Ѹ�%�됻�E3�V�iB��V��$>{>О���N������N{O`YKe(Z����G0e,(�g�A��Q5�e/��E^�7rӼ��ꉌd7�$�">��� [ع����k;�=��C���$<=�:�r�R �ea���ě4e:�Js[>�@��Ѕ(���7q�C|�4�Q�d�8�B��~!PB�UMM�@�Nb�S�qW�։�ᢆp�"F�|-�ҋ����t�{|�z�����2S=Sz��:��d=5�|��D�G�`����E��w�'�`�܋p]�=�zG��y�|�5�>R�筩�d���Ĥj�K\����R��O�U	 �������`����(�Oƛ�}��+��ҴVe���
�K|�}���/x&��8�-�|��T@�G����K�.B��Jh^8�r�RI���=�	�g��7�$��4�<�Z�XM|�
6%>	�S<j�ea��Ps�1'R͡�o=~�z�^�&�8�f�.�"6l�3��}l��A�^���̕?�'1j,��]��fi�)��b�+'��$�'�hK�G��4ښ���ҙQyR[�P�_��M���0�,�DH�`1N]܊Gn�Ƶ+��e{��<����~�.�,4x�F���`�� ��i����j���W�q]z-�OGb�;�K�}�Gí-����hJ�Om��p�����~���qbw'�PK"�J��Z�E��겂1?���,���T�#}�h(�s�Жd�:��!����p�C�Ƀ�"63�P�c���zV0�Y��0�	��z=�=-�joC-X��lo�
���H�qZA�6�C�LE(�4��@kN�=<D���,Ź���n�&B�p}��	ΛD�mb���6\�ل���8��
'��C%�=T���<l���(D=�h�ACf j��դx�!��A�-Eo~0z��~�Y��/	�HUFk�0T����h���9�Fn6�q���;�I�v���yΑ�g���!(����<n}���ߖ߽IA �������`M��y�4~�/?�k�>�����k�а{6�Ag"�I!t4+��R�l8+GR��!��lswN�;����������ǖ��Ѵ5�P~p
��#zS̫�>ۋ�Ǳ����q��~���4���x���`��.���b4kg�@���=����8��-�x�i<��8��U�̴��#�o�q�_�R ].��y���d�E�D�(Y�w�z���R��w��K ��`s��P�� � �Y�r���r��Aڶtn��~�sMS;(hS�~.�T���$5���S��sp���3̟8���s,��G��>��\b��&��K(i����+�?��\9�m+�jiV��MlJ��N�<�raZ�Isg��Z� J|J�)�֖B�#L��&�c����Y) JQ]9�c�?+	QMS\�]ݵtM{��%�:t�܎�1kj#�Jj@Yf|�,+Xn\+Moy^ӫ��a},�j�a���D�i�/�rq��.���x��'p��	����8^Հ
@͋B`Y
��%Z�D4C%*�[�sz\uB�qiUG�}5(�S���2dq�܏����4��*��-ǃ:`���X�h~9@;!��?��a`l m#���Q ����d�-Ԁv�5�{;�B\���U�>�Q�@kAe(�Z����� Z4	Q�S�)��j����`����:܁�c�h9;HtNc�K �uqP���:���`��	�����w���W.`�s�1qc+/oT �f����&gF�t�y�VtS��1~e+�{Ka`���$l;������}8s�:�ݺ���ɋ718���[@gv���g1�y/�Z���^J|� 9��ō(��@Yu#��S������m{���4���od=C�jk��܄���4�cfj
�/]İܦ%/gN���/�����`hx;f����s��W?��?���+�����!����x㝯����(MGTl��jT�fV^=2��Wڊܒ6�qi���ѤB��"0$Y��[�8���*>>iY�(.oEfn5�s*02���<��'O�erB�7-��~��q����Mt�Nw��]kl9�G�;��K�q��s8��l}b�n�w:��{b�Ѕk>?�s	�vI�A�C�����9Fxr;/ �m�����l�y,o�F��F��-h:ҡ��JZ���~�.i�{�(%@�W�BwYkU�+��^�ƒT��[�)Mq	P�尘�9��`�>3�L��q��?w<G"̊�4!8��Pm"T �v�k�8\��>�����@�Sj@9_�D�.F�]�,V�	Jo�P�>�������PT!e�7*��Ý!5�w.��,��yTK� +U���oI�Z�Mj5	PA�'_Ë�۪�j�e��#wWn�� �-P�j� ���-��	KA���5�XPwr���#�$n|N�0��S"���@��Q�HW��8AȂ�4��&�ID#��O��7�0!4=c��8��a_��7Q�x.�2w��5��R��E�zq�;�ypڛ���$�����":������PUJ�rzq�������@1� ��3�	��W2���	�8�3�6��'{��O�to�&�`-a)�\l����fx�y ��T��@J��	��6�==0F�L��`�D����f���0��Ѽ7�2�NԘ �4�eR9Nt�J��,����5R��k�x[��8���aD����|~�\$6��|�
�[�ۓ� �h�f���� '�m�#�ĥsh�B]�m���\O��{å�ΥAp(�]�qYX�7���0��O�چW�؍g��ԕ�$4�Hl��gG*ܥS	ԝ.����K[p��6\;?��<��i��HP����4GuF &�qa�gjpr8{Z�1���K�F[����F��>�D��h�Eh)����n����dB|m���������a��^�(�Ge�:���
|��`��;�p�/����
pz��y�0]�����F��Պ;���f�b���V�ܶ��Z���80Q��CDhg����_���0t�+xvqؙ�n�'ӑ�N���:��������b��:#�<��=-�n�s]�ٙ�ӕ�k8zZ�ş���7�AQ����1�wg�Y�("@㰆�o��$�)	�Qn v�9�_��W�����c�Ž(�n�MS��ځ$U��9��F����U��mL��'�ޯ~���~�e|�g������_�	?����G�=��Ɠ?��G�#��K�����?����x�/��ﾋ~�>�o����@*�����"��#ts=>�౯����6N�y���aҖ���o�R U�Y"K@Q��ZA�ҵ�+��^������o�Y
�� U��2�MqUSP���C˝�p�\��=H�þ�'�O��G�L3��O_������L��bCbU�+�C��p���ѿ}�gw#��4��w�aW��5@w_-�vU@gg%����X������V�����q�D��m+$Xy,,D�9&VNe���t�Ң���@T��{7éDh*VI�c�
��FW�&a5!* ]%�q�bԵ�kZb��%k���X]�U��XVr�:�Q���� :��A����Q���q�cx�'q�8L�V��#?va�(U�p-
Ba�s�Հ
@s&�Q6ۨ �j@����x+J�עhw��h&1���!׃&Od �?a1����.��-V�A��j�
��~l�� �&@�O#C��b��생YV�@TE�Bh�����(���7���8Ay��p�ZM@�tq\��vl�RU5���B(#����z>N�Y}�S��� @��� =7��u�ڴ�ޗ����gx>&B�?���R�)5�����*��:�c�#s���^�l�˃i���E�83>���߾3g�i�~�>zN^¦�#��G��,'����IY�HϯAec�GQ�2H�"��.�pp�FyM&7m�Ԗm��w�Ԥn�R�ڂʚ*t�����V]:�u+6Mm@vz�����㷿�G��ګ8~�Bj��/�9���������m��hnnš#ǰw�!L��m=����[��mAG��KZ��fԷ�����i�e��I)ENA�*;��_��ԍƖa����,�m؉q&��I�ؼc/n>�<�<���^Ė�7=��>��v���t���Z{��\$e�Cw�����-8��˸��m�=����F�_#<�n�+-�/����i��au���]�t3����h�ۏ�M�g��e�E���oF��v���4	g�O��Z�n���@���}XVW쏆� �1�Y�
�E,�����z![��BxJ��#ma�x�x@�	�|-�@������Mz�z�"B�I�ۻ1�:��Zn���Z��س�q7C��L5}u��g�-<�;7"Ѕ�T�$�<8_�y��D��E���B���\��q����FF�)��M>�̗�M���~Js����'C��iU�f(!+(�ҴV��B�D�ɴ������Ni�+���~:)�J�����O�>�/�>R3�q�`s�2�ZP�ɖU(e���{��F\�+LJ��`�E *]"���+�E|����k2��w7^ħ�� <�	O�x��yhjF�j�+Mu��.�A)���uM�&@�.��w�5��Dw�r_����!q�6��B��p��� >�?���F�<K�������lE��C���>��P[X��<LS���M��x&9C?�	z�O�#�	ӅȺF�DgK��8G�:���#<u����`�� � ���2��|.�l_d�M[[P5RJ\F!�?ܑ����Ǳ3S��ҙ�ذ�i垈(qG@�?���L�:dv� ԕ�t��D�[I�6��C#x��&\==��|$d��.��_C�Ѐ�l���y�H��Ƕ#C���n\yhíɈ�և��r�X���b��?U��؆*B�����1�8�@Zj��PKT��w7A��jD=�p�e�&`B�`�d��|5�y�&��a�pu0���jX����J��"��s���h[4q[��yc��w{}v7'�`g:�����HN���x1�N��!�6t[���}�x�'�'������ߎk��>�84^��E88V���,]9�ޑ���,lnH�pY��fW^�J{�?�3|А�6��0=�Qh�E��x�"�m�u�.��p�4���1�\,��n	W_9w�  �!a��½H�z�v�qe��
,\��bY�̋ñ��3��~�����[�������;3�����,�d�4�e�9��HX���x����s��*��u���W��w>Ʒ�#������?�W�=���o��#�q�H��W?��?�>����x���o����_Eˉ��X�M�0�Z�e��t]w"b�[q����w��S����B��^��gCk2G��n/Q���w��-5?ҋ�\�(Y���bVR�&�Q �<��Q�@rك\O� �lA���/H��s\￐��|���B��Ո.֊
B?��6�'���O�sQ�b��rAì�Y��;K�zW)Vn�̓�5�ʰ��+���;��!k����Hd�ߡ��r쬀��Xm�B�����B�h�}�U�<Uj
�z���Qh�I����,�o��$�N�OӉ�)׃�˿������/1{t/6>��gg4���U�����X��R!T��\?����j����r1�5sD'�k�8 R�#(��y�r!�6qzC&�Of�X�������X��ʅ�Pi����N�V�k!J��YD(��5��ڎxU�v���x� >WT�2XU�5�nM4�`Ҙ �X�ƨ&�6E��.��G╯=�;/?��Ϣ����KQ����Ӭ0�<oe�BWZez��"~5q�K@DSR��=V���`�x��f4=ԃ�ӝ�<҄�=�|	���r�#{��SوLDDg,"Z���W�N��	�\*��^p���5���++5��2��S��� TƦ�025�z-h�h:!�OQ׀&4g"�3����z���QMp����El*p�N���vޝ'5���VSS���ZO�V�L"��
<����̀���͍��M�4ץ��ȸ2�:n�<r�	n�iB���c׷`�sq��s8��YլS:'�
65��r'0pqRݒE2~s[��F��q�e��-�m�=ش{��������6�o���ç���aϑ����Q��t�����m
�c(��Q(��Pi~�����Z�s�����@�S�-%0˫+�DT�r|jr���FKS�==0;����_������'ٿI1��C'O�_~�;���?@o?����FO���k04���E��fl�ه���HϩAym/��7��m��w٥HȬR����mF9¢2����
J�s���)D�f������]��ݻP��A���-!V�n��#m�^Vj=��@Vc6.�~;��Ŗ�;p�Gp��Ә�=�������c���X�yD�!t���_���ZO��Ch��b������}<)�d�j �ux�͚۰�����)5ޭm;ه�������X'����*��C�W Z��:!���Ey�
ҽ��BwV��\��$��ln��PDr��A�(MpM]ta�w�%*5�j�����R˹p��`>�
��A���}Ğ���cBו�2�=�F-�`<���d��B.<V�]|�ĉ��K��Ԅ�U-���R��&�N�<�M ��n���mV�7F�	@�\.b�;̕�ՠT���ar���X��A(��y��{�]̽׃.vB$�u��{Ï�>1��t�a�!�J'F�^j�����j5�k��� ԃ��:����D����$�QbT�ݺȼO��w��2���ħK��ZOs�vTat���o�?|���p�W:!�P�xF��r(��|r������W���d�G��ħ$� ��ZaU�%օXB���A�%�hJ�Z�x�4� �GiB��I���0�	�彑ZP=��B���:D��?�{U�Gl�FYA'�z�a�̸�2Ɓ��-���p�u壠=q呈,	�v�@QC"����q��(�7� ���6.�G��r<����� P�ԫH�S�L&6���ʩA<qe
7�Ʊ$� � ����wG
�?Թ0�U�8vm�1����vPg��p4[Gӕ��BV�#��S��F\�m��\�Յc,��	V
���(�v/�4E��z$��B�쨧 ��cA �j�73x �nfpw�����W�R9\M� ������<�uܾ�����Tq �VF�I8؝��|G�cC��x	NM��iB�zЧ���9n�����C]�����u8=]����qn�
�T��D��b_o>��eb�.�� �M�凖l�����Š�,�9a��1�Kl�3�x���9��N���1���	j/~�����AD��(_��|c�c�,�:5Q�n��A[2���m]���_|��>}� |_���1|aZE�XQ��co�jv�l$	�ƒ���,��m��e},f�8��������Go���_Ó�?�g^{Ͽ�"�{�����x��W��+����_ŭW���/=���~O}�&���h:��m��#�M�0�� T��m.�^b�_�x����u�гo=��]}��Ʉ�6M3D$X/T׽-���{�\����ij�d��r��@A���A�a�:
}
~D�}��Te	�.��W��I@����t�- U��*�Q�Y�yd�G�Ѕ�;ˠC���l)������Y���׾�)i�i��j;���bB�F���,�o����܋O�����O�g�|���?���kص	�摴�s���CT��l�� %�@o�sO�<A�L�"J�s�E�ދ��SYXN����,r����BV�sM��f��55���PA�"@;��x�w��(R���R����P�#�Q}��ǰc�s�5�U����r�4����y�����ƻ�U{�TՂ�B������'�}#@C�ٔ���|�N� ��Qt������� ���F��2��\�g��!mc�FR՛���8�x���k@�' �#�ODz�N�2�O�&vf�z�GE������j��$0�^��#�b�ۻ=�. U�@��Szo���·��'z��¾tB4xki�v]T5^}W��v�M'��N�[�l�=��®�`��}�Ɠ��,��G2��_�R�{�ʽCǯ�`��&�T��5��5�}���>������o�s|
�fp�����%Uө:J.@jn��PT�A�v!��NՈf�W�������@aY5�<�����T�����Gi�+/U �hoř�'q��~DF�����?��㿪c�����MO#?#�9��02�cb��C�C8y�48��Zdd�cxd���p=�[��5���z��F��������FFQ+"�����$�gU��R��_܄2~����!Q|r!�6���k���lܻ�M��Og96�,����H�j����˰�b-64��[�0��n�x� ��	x�Ư�h��zE:��X�f�E"��g��t^�>�p-�Ԁv�P�T:!���~��ܡ���؄��y��! �F�n�֡jW*w5���9h�.U��}�S]:��� Z�BiM�j�QM��dx���A֔x'$���Bp\��Y0�D(�!���f��"#����X� P�HuBD���$B�zPgP+iVhg�������
����4e�#6	E?B��JE���,s�����������$n'.S ��JM����r��e|��Ñ���G�������7B���"�tc�Y�)�o-�=��\@������@TL�T��
*��ޛE�J�^�D)��HD;�O�8r�P�]È�pg�E��,�S�3��@8,�1�	N��p�/�Q\����Yǅ0��t�C4�źi���ӌs��*���DP�p-�[�7\	O�D"3�VQ���qV�o��:M��kA��aA,�s]O��#.���"4�����Hs,���|+"� ���=� �/���V0	&@c\`��s>�I�+L]`��#B҈Ǉ����՗��0�Y��ߟAi�q[2|/Fְ�s:�N|M����3?g,S�_���x�T�"8�9eؿ����0A<&f��?����.�[�/�
}	P8r�{E�	τjB�.
[w4���a<}m���HR��Z���P8�u����nJ�gy8RY �yjϼtW��DG�$��v��b�N���n�q^�h�á�*\�����"l�k�亣5њ 5FY�	�,P�m�,{$[�A��2���@��%A� ��}�_������>������|=+�U�3Z	o���缂PT����"�2<0Y�ٚ�iK�"t?s�/�F
ql�'&Jq�'�3D�e�Po�h������7w6��l-�o�Pײ��.�٩2\�����"����,��4L#�fOA�hS����]��dU%��85!�&"S���� Gx8��d��ā�����.�1�@X���?�N<��D��<��u��n��Q��!����������m<�޳���c(�i#@��%�	�Q�ut��iX1��hK��G������}�����x�����׿���{�~�^��-�L����}�]<���x�W�������b��!��@ĆZ8��zcL�˰b:Z, 걠h����و�҈�/^�ӟ���?}����a١�h��	HՙΦ\�ٜ�� ��GW�����X����=
P
��4Y�?ҴU�'�ӄ��|X�_���)Y
�*r��gy���6���=.����U�\���w��]&��ʼP�gY����J-�֮rSF�Jᾫ9GGP6׋MǶ�g��Kų���q|1���"��Od�K�' ]�� ��r]������zh'
�#p�6;ja��� ��P-t-�F �}�����Ⱦ.MΥ�f��y���{�|c�B�
Ɇ,�\��	]�j	�n�"]@�j�+��}LO��k��uD�tF��P�/�j��&
�+#U'DPú8X����5�%����EHW�����f�����mX�<|m������ u�My���4' z�n0`�J�P'� MV�a��k@�������h:ߋ��(?҈��5(���Y�<�(�k�I��gL�Ʉ[�7�[�R ]�����P��K�;�K�4�#���T�փ,��5�D�@S�zr�n��mY�\�"B��"B%�&��Z���O�g��>�>4��� �ݗ��wu\5��6�m'��N�=4���[���l~tq)���
�*	�����~5=��k3���UZ����h�p/��6�|�u\x�	t�9�ݼ����gR!3<.���6,r;O�(CdbR�ˑ��������m]x�g�c��v��N�$RZY[���475`vv+::����G;������Kx�Σx���yt�eE��hE{c=�2�\׀�����׿�{�|�����䡵�۾s���(��B^i3��j�ETf�4���u]�^�J�$���6�
�=�P���~�Q��r+�W`:��(�:�}�Oct�,
�����؅z�,3��+������f���W�{�Ѓ���o����a��f\�P ����F��] zylai��@��3q��A�����q�w��n��>s|z�n@��Q��D�z�M��_���-�	n�fP��b�V�m�	O��~��mXjr}P�#�y"7�Y�p�v<�1,<��m�aX��Y�5�_�ae	;_�����]z�z����:�����zp���5���m4S �%P���6[��:���$����Yq�죁��LGƎ���0��B�<M�<���^�
��L�=�2��K��ks���B._���`��sq������V�;�j�I�(A" %�|8�_ J(r�5�x�'9ω�Y���v
�r����u���6���0��?����
:%���g�#�ehh�^��/�;X^�V�9|!�N�,_�]����`�u��4!Hm#�#��Qΰ�&t�����V"��
F�R�*(u�s�S��en�!>�P��S��
>;!2�# #l�EX�'@׆��Xi�jA�DY`e��|Za���V5��ċ%�.5%F-���a���u��8��?�A� Ӟ���HBpE��8�F�60
cB����i�2��o����
G��1���q�\���D6�%�H+�F}k��c����~l�AV�3³	�Bo����$΅~�	�m����T���d���Gx{��f�8=�M|��
_ԓ �Cu8k"�C���! ��R�����R��ds��9����[���,G����m0U��K3-87QNF(��%٨�#������<$[�E�у�_�([m�8!-�	I�hl�3��aN��yÇ�qq6����M���x5mt���8�	��ߚ�_t'�`PZ����s�lMƾ����|b���s��'�N�����������$�:��C��85X����ސ���Xl���hY8��Cё�6B��,C5	�b���<-��N'@�����@wz:��ɖ���9G{��!2�Q1�<��!2�QL���|�V��Ы��vs<;S��<f�/��:����S|�g��ŏ_����ޞ�����9$�~
B��,ߐ��]�ˆ8L?|����x��o���^ ,� B����y��w��?�_������}���kx� }���������'o�h�V�Q0o���JX���	�I�e3�Y	��2Xm(D��n{�^�6���_����F��!�I�b"UoG��Rs) ��&���S"��T]@�\�(��G�B��(2Rø����es�K�(����x�~_��r��R��S�>W
2�=�§
�)YI(�$4W�^ (# ]�����m��Py^��Q/�pM��x�e��P��g��UL��2������E����R��Z�^��'�|o���(����/�������>8��X�T�`G�w}����Jm��Y@�V��3�P� ]D� t�t6V���S���Lfݍ�<�B���۳��wkB����g��IXם-IW"ַ�c�ⵠLmVWi *����gޢ�5*�S}"º���B���xϾ��ݹL�ë ���-�tDd��� h'�@/�E5�iJAhC��������zG��w��F4]�CZ& =P��}5(�S�n_���y"ucR&s�:�O�n�X��mX�' �₰�h$�g"�)C�~g�OM��h�<��w�§�R�Y�����v��mW�Mp5�-�W���m���h;1�����=٫z��r���c�9��* m�c:N�'���}D�8F�l���-
����о�
�Ϟs#*R������q��OZ(L�m0wt/^����z� ���<4���bmXᳵg������a�J��f4v�)���U+�Ƨd#6)���2��o�����46�&���ݨ��SMp�2�P\\�Ҳ�q����u��GlDRcbQ�����bԕ���	m�(�����W��?�X���o�[7�Dc]'������|�q4w�!1�ɹ�(��BBVB��׀ȴ
x���=V�>�%4�J[T�grZ)��<�F��}ϼ�^|��8z�#�Ȭ�@Pv"�0OX��A�R��Wb��ep�����n�������{�<�|��>��k[0rm#�	~G���(�)��� �e=h��5�]\. �f�mG{�mX�����٫n�"Mp�O�ch?0��=��6,�n�|=���TZ�5����@B�慴K��Tn�R���4$;#=�1��tr��{p�����B|P�9��O�@C�����g/��D���!t|>Pw�!�y�k@�"=W}u��?!ɡt2d�KW]b��yI�(�I�ۺ�n��sh�ik#X93.ưp6���,�a���nĨ;q�!8��6����ZG���e���?�e1s����|�'s'#+WS�3��s}�7s.���ĺ�%���-+�GK7c��9d�݄��\2�NY.�#�	S�}�&�ְ�v��1W�qkح��`��W_��Z�y�8mJTޟ0�S0Jt��J���mK8��2�I�)���Ԛ�j�k �@#5��QD�Ԍ��1�p��P���u�-��@{�aV�&�­��Y'5��VX!Mq-�Bj?���S� 4�$<#�`��ܖf��|�V� �,����	�iChF;��2$,�@�4���I���Cma.ۉ(3�&r�`�YB?���0	� K��lC�`���!�N�'�(1�>L�^�R���֕�}��q��8n�cK9�˼�l�|/u�"?8�y�6߇ ��#�S��/��yarS%����wb~��m1.p�GE k��\��x��Z���LLo��`w*j��C����Ձ��\���k�f�Μ`����ũj�j��X�'ړ�V+�(�5@����	����v�H&<��@B3��V:�� *��X�����y���DՈ:Yj��d���#���\�,�����HpBg�#z�]1�㋩�0l���|c"�tf`wW&vr��3{�3p�?�Y`���ɱB�bN����@6���@W*�6'b{M���X`���;dT�C�� �9֘���T���,��)�ȉ�AJ��B�����o7W�x�!�<�!,�]_D�#!)1	a��K,����i ��>�㰢$V�8��%��?�O~�C|�g���WCֆ:հ�؛��}�X6�,ր��+[�`���+��.��?�����^~�o���+���	�=v��=���_������＂W�o�>^��M}�jNl��`>�3a2S=F�������L!�u�bYMB&*q�ūx�;_�;?��?zE����4k�24���*W5�r-����_ �D5�%��B�b�ջ!��ç�.���>ǒ��[r<�� J|��k7��K T��й�k�U(��y� �?ʗTw%,���C](=>���^���Wh��"�d�/Y�O�}y�'�Կ��[
�*����٤�����_p��G0}b'Z�mF܎N��T�dw-twWC�ǀ6�}?@�>��s�*2�ZAT��/v�u/@�O��E�Jf�D ���\�j	*�i����5��T�!B��r�^�M�vo
�����I���c�ܒ��������� �N��	�]G���ٖ���\d�`��F<��x���wk@�J�\ۊ(��4�5ctx��It�0�pf�>�Y�%
���6b���.j ZJ��C	S,�]�����"}s>2���bx�`����9��kA�JWՀ��:EՀƷg�j��gX`'�>��'��cw��
4�U�ZTm�\*8�N���;�@{�� t'F������4�D�_zh/�P���d7�w�k@;NI�j��6l���K|�%�0�97��y>^B��12>D�L�چ�w�aӹ��l.���-������`����B:�ym� �x�����ٛ�x���n@V�4k�GNI#
+ۑWւČb��w��?�����Mh��Ce]��H *��/.Blt��3��ڄ�s8~��\����$Ų�����hT�䠦4�%h���x	^|�Y�Ɵ~�<r�I�M��gc�[QQׅ�n߶!�����h�DzQ#"SK�X�R�1�ۏ����$�##�%m��m?O��V��<���n����|���{��z[����:F��������:��[�ek�!�*/|�5�}�
�>�g?����^ƶ'�a��f�^�V �k|��ݽ�����q]�.����,��e7f�Z{�<��SS�:4���D��Q4��C�U* m8 ��܏�(�J��]��L)Y�]%!h��Gc�jR�P��0Ku�gh0���X ,��q��u��\�iLL��4�6�����z^z���tB��m]�S[�I\���4��vւ����,�bW)d�ZX}m�ڮ��gJ왰pil�#lehl��q]5_b�iCN��8߃�,�#�	P�~��BB�Ŕ����F#;��9���xc{��D�|gLױ���e�>!*�/��&.����z.y���g�}����=ibh��3��k�`�Ϩ���|��D����K�Z��[Ɔ����dܒ7r�g �M�iS��\7G�[y��&\�Y�7��Z��p�"���Z5�g�����e\�Ys�C�=�aH|pc-!ԬTl`�i~����Њ߯%e�q5$�dh�8�����"�~�DJ�#�4��%���B�HW�G��.�&Z�	U�`+�[B'��0kh��`&4�K�ﮋ�!F�O�~.�E��"�`&��f��0#ح���V|�愣%�mMTK4���#.-��"Fƭ�9/�Ϸ�p�9�˖�㶱����?p���k���s����)�}LTk i���q/~�ԼPt��g�U����J�ܦR���ٽ�p��gKQZC����=��p&�M�o8���< ���pK�Fp�&X8�~~Oݘ����l,@]g<3�Vw��.��km4<�B�C�Dv��E/E)n�#@�	h���ׂ����� �A���/MW���3��Q��A}�
|��𢡊� sT���4E��>b��`"4�z=R�,���PWd��>��vVk��󄷻��5�������|�x|%xZ�(�M)!h��Dc�;�Ѧx7�d�a� S��Z���$U+:ߔ��m��ّ�=��^"{_O&�e�@o�w�cO{
v�&aWKv�'aCQ&
ð�<���*�Di����D7�c�9�!ȊrGF�����0 -@ҿ�y#��A^�����^�40�^ގ	�B|l�b����X/Xd�È�4ݶ$�i��jWV���>�z�|�-|��q��H*�AE(t�c��?�$�I�	M B��~*����G���v|��O������8|�8���a��ݨ<zULq ���Yhو;�����x�;��_� ������y���2��'[�a��fEXV��e����BtG)毟�#ￄ���ν�$jv���8J���h"W]g�
�D��)�J�,�4���PA����A��D )�\�^N�-�{�R�j;U��d�Md���.�G��ϱ����洌�w%ד��RY�B�
�)C�����k;��,VY��X$>�Bj??7]�9���[��*���Q˘5
����wO{*�ǘ﯁�rı�Qyhms���O�)4#È���d\�-FS�A��mQ|�w��{#���?�U���ӿ�o�f��b�m;��:ậ�c��S�]U��Y��О/S����e�����ܮH��u;J���ߏ���y�u%�+�p�!��˭W�r�nc>�7����,��MyX�� �%�N:�bt���.�Ě�t�΄� ����g*��:�)0�I�~w*���4�'a]]��EC�!:��e�aќ��d8֧ ��I�5H�Ė�[���wp���C��W���X�U��,?z�>0���n��C��hNEtk*2�
P���]n�>����:����8܄����z�E>��M�gϖ k[1�6#g�<O��\�u��5��^O�
,Y�'.��O�L/�ST��p�܆E�ilfCmh[j������xDU'!�%�Mɨ�o��I��U��]'��|�RzP���]��ہZ��@�Z�tX��>ۏ��M����ڸ����� =>��#]�c������~{3��N��rMz<�tB�wU�"�����X�0���|���~�'0����	U����#�72��|gv>q�s�e9,"/�/�ĵg�¦��1�e;�v�Ц�jDu�0����]G."��)�5��V��S��"��I&��}PXZ�7����x%�5��oAS��؊��V�����O����C�74�Cǎ⍷�Ƌ/��C{������h(�DMY!��1�Ӊ��,���+�ob����1�u���a��V��6���9EMv����mch�GJN�������
<��[����=���<����i4u�br�:y���Ǚ�����1{�0Z'���T���؇��E���cs�6^���a��j4����O���N�^��~�1\��c���>~��6��s�����x
>��b�r��+�^U/�rK�Wg���u�'�6B��vk;v?�#ܗ{�M����s�;8��m�w����PM�������Cm*��1��6�]�=���G�š�+Fg��=��ମ�������PK�ƻ %�q�^�q�G�9�=�aN|�y���1c�yz��qc���MxJ��:gmh9���������Q���pgaܝ�p"z�<͸�PG>��6��5ѻ':��U���uy�'<}:Z��V���k ���@'��#
u-�#�6�y:�i=+=�rB��jp}�ӳ�:�|}�TZrq�s�k�3��J#�Ky�����֫h/.�^x.�{�����]bҎ�gK��&����06w0TC�6�g�Y���FGmCA���rGBԉ�'�{Ƙ����d��|�a�Ktz[�ȴ�֛�$^{����r+"�Ɨ��	)�Z�;bՒ��9��X-L[�L�� �R%W̓�e���S�#�"�����#���>�@�`Bx�V��^���=������c�C9f=F7\=I�	T�H�1ډ�{"7�	�|"с�v"t�{"�mb���P�'Pe�D���wk�%īU ?��BK6?��B�k��X�y��cgo��^Fp�1���	|y�y��7�����zu^z�N�J��OW�|���,n�L�	�!ٖp��O�:���^p(�"@��R��Rox��"���;�q��n�G�Oc#��,�{?׷%@�PԳ<�U1����t�*cQ���$W�G� �U�i'MqW �a=���74f��XvwbsUF�C��� C�!���v+�~��j�;���D��r���"�����C\��� wsxr�r6B �G_wSx����H�Y^(�@ӐD��1���^hN�FK�':R<0�s�$;�*±�*ۈЭ��mr[�y"u��2�oL��ј(��dE�8�c���1Nt�4e��<�,h�' +�y��(ɌFNR8�B���� ?D�#��ADhH����3$�����tL�?�"���	�/؂`P���Xݙ����ml�F��~������o���~�]�}��7���"z�1Xן��IxP :��e#	X=��խ�0i������?|�������gc;�Ϲ,�AwL7d�x��҆x����[�⣿�/��c<�����g����z��v��5:��̇�X	t*c�<ߋ��.��G���o��'��������8��U\��%4]��~s<tF2���ph_R0�"@�P��"&�� Q�yPj���F�G"vG�ʃÿ%��^�G�SP�@����K��j2�ɽ �7�l��|>H|J��+�����Qˉ�U���}�
5�j��<���Z��{� Uwᴧ�{�`y���*�z�U�X��9�_��ϤG�}>´����o�_�s���������w� ���"s��;[a��F�k���RE�#1*׆�6��hw5�S�К/U�o�t�<Q*��)&(��o*��-�3n	�Xڛ���"hM@kct����VF�J�]E������\���ڱl����	O��t��f@{ �����ˀ~W��r`֛�.B�=��I
�:U�Lt�5=�Z�J�'Z͂4�y!mH�E|k!�O�≯<����¥'.ct�B�R�R��8ؖ�â0
����K�v�Y&nLAT[:�;ґ��Q��Dچ+�0~mZ5l8Յ�#D�^t_�hQ�='�)�fq[�MV"�(�-V�m�t���P-s���t�]t~.� �� Ԅ �5bِeR��W� �1��i��oC���=�	m��.�����n8ԋz�'�)�%Be(�$����� <��|l�BZ������&O��Ch<����n��� Q( �=�jA{ ڵP:pm#����9L?9�ч7���l?;����K迼�!l�7�p��N��1�g����p|��y�}�(�NOp;��;5�3c8x�!l�w�3;11��vE���w��
-���_Յ��jĦ3D]&��󑐞E�z!26�<�2�<�4*��PQQ��vt�����)�i�(��ǟ|,g���k�/.�������������O������y��-EUiz�[��X���
|��R'�_��W���~�?�x��瑕S���zd�7"9�
���ކ��z�d�#9�yU�w������7�D~E�c�����.��w��k����;�?��s�sf�=-H�.BPF�b��r�'�z��Xn�˴���}� ���:�j=/}��}�6=����������iZ{/6��F?7_ ��c��!@�q�#B�OKM� �8�m7���}�<�}��	����@�:!���r��:P�Pg�����D�~��,����ò������pY��BБ��u땔ıP�zr�;22����p�'Ȃ�fCX{��cN|�y��	�i ��tу�;�ClZp���t6�xHA����
��;1�L�8
=,`ZKX��ĒX3��|>WUK(��P����z5m�j� ���7қ�eI�i�*�H����<]+��f��i]��'��<��K�	C{O�m��.p��h,5��Z�R۹D�̀�K������Q�<�Φ1���ܦ�\5�]i�+��f���x���ń�������<�nj{r[ʶ�%:�l����Q��g�N湰��F�u2_����2.�������c���� �P�E�rږ߫�Km�԰ZZ�R��jR���O����D��>�@�A�p�vt�=ߧ=ߣ#ߣ�����P	w�]�*MikQ�봊p�%ai��pXp�2ʙq�5�i㢮-�kM�c9�N��<.�s��B�-8�霉��m&̈́G���s�\�I���y�`TP*����&�y��(�ʇ��{������5�+������^Dh`���b��9>�k�qp{#�V���Z���ɹ�^�(��Dx������\���<O�KMh�Ԇ�£���H,���]�z~�����6l�F|�#���R�OԄá>.u��@la00�������0K%�!��$���NoG�0۬E �a.��I��\g���a�8�*�Eo�b�PF|J-h1�^�g�\i��f�h��
�ak�c>��p������3���t2�'��O��{["�Äw����,-y�>��'B�C��`�'��:�U��k��7�9�=���Ĩ/&�É�L�p��&��t�$���5��\+��Di,F��џ���pt䆣�Ӄ5ik�� �]W��d?�&0��|_��ȉG~J$��=��s�� ���^�pCH�P��P0�拠H�Hy�*����0l��P]��h��iY6]܍o���ޏ>���|G�8��Ip��-�� t"�'k :����QЪC���x� ��7��?|3W�£)�,�Z�0k�� &,��&ä;9��q��gp��Wq��'�ȫO�鯼�O��x���!}k��Us=��<��O�C�	��_�O�3>��x��q婇q�����_������o݄CW&t{R`0[��;X �g��#i��r�M���C�-��Z��GSKzo�Q��hj5�F�Ryp��X��E(��s �&�� *�[S� Z��]����i�UX�h�+�����{k`�� �_��5H;ٍ�]�7�?������ �����z߿��?���S=:��������u0tK�{j�M$�l�����;�ѩK<�Nncv�\_�(]�U�Y��*�n+Wљ)#,���#@��K���X�R�p�vK!�>7B{�8���ډhs����fB�7�}Y0�ɂ� �/��90%���Ӱ�*k�#��r�VA(V��bY���:c9˅�3|��}��yN�$�B���:T��jl95�?~O���=s��㈭ˁwE2lKb`QE�JGD|�TP�M\h�Crw&���a��<v=���X�C�C��=ގ"n�n'
@s�KgD
�Т�G�3����zh�h���m�V����6�"�"!��h�ۇ�K��utm��t��o � S�N��\�g�^��}b� ��� ���c=h>ޫ �{e������9���c�{��}@��8q:��n�~�6�ي�+�}~L�|4�l^݀��,�=����@�ŧ<v���}�v?ye�</�w6�:�s[ �ݰ}/�Ƿ`��޺�UMO)@r^�����W���\��e $:���Fz^B�������>�_��kh��BYY���҆*b/;3c�x啗�����s=]��أ��w��g�}�uM�K�EYv1J�
�P]���&d��`f�&��R'��_z��Ώ����AL\b�J��Y�Ĵ
��b���HͪDRF)Ӌ��Z�[�=��n�����9E�
�Y�u(�nG{�����z�-L�ڍ��>�T#� ��,;� $=v~NXc��V`��*��W��7��ѷ.�[��z����Ob�m��� �B����\��9�A�yA� J��]G�0s}�>�c��S���@�\
7W�۰H/������_
����
�G��N���� t�"�<����љ�r�P
S<�Xu��$wd�z#9��<�G�#8�����w�5<��~�ұ�t�c�)��,��X���}���˂������o�C�3��D�W����	w�7�݃�4��,t������,]�Si�J�Y��>v|�������)�g�B�Is\i�*�X��T�i�g�J�9���C;ο7���p��{�s��q�qG/�I���8xZ�y���pca��h:'�{�j>�g����2�s���*�[jp5���Djt%�|.�?�����]���2O����
��O�������ח�����
%�8�7�万Z&��|�_�'<���Sς�[���?�t����:l�U�0���'��8��3�q���2^Q\7����y�\�+��'�^�{��"��Qr���	�+��	,��q�1|��g�7<���W�%���{�9�C�E�M�����g��z����61�#/�/���}�v3����rS�Ռ��T=W,��h7uk7Ɠ��[n����'�v�#@}Bl�d� �������1���1£l〨h;�Gvu���Q��ӆ�;jqqO.����{|w&'��W扠4K8��Ds�+�s=`���<78�+���L�m��u���87�sǺ0�!љ�����
�]]���Z���&WF����5񈋰F��!2c쑟䊄+����E~Nz�!@�,�#��=e��7\�C,���,�ֺ��35���(�@��%
��CH&:�+|��B�����e�� gd��!��/������x����}}-d��x����(-e���NFCj8SCQ�� ڐ��:~G��.��rbК쁎4o��`�0�Q*c���f8��~�s��<}��ʉ@{v8�
c1\���,�V���4u�W�'לD���KDAR(�#��CC��y�"ԛ��ǓC/��z! ��A���El�?������s�3��aM$�Z�ݙ���Xߓ���0*�֛���~����{�}{>��lԄA�3k��ħ�T��6fbm_<VT"g/>�������c����1��x��°+:r���,�;zۈ��w�#`�����x��W��w�����S����S�qIH�@�X-^������O�7?yW���Y�W�ţ/<��~O��"���޺��=�Пʃ��r�H5ŕ�Pթ!&���*\v?>��K �>�R�p.�s�BU�X"�^������HM��u��e}�}���/F-_x��5�+@%j=(� �y���*h�'x�UB����_�5�8P��u�8݋��ݘ<:�o�_��ot����q��yl9w U�.~�-�����-0".���A�x4�)��;W�-e0�B�n���d	V�g`�p�6q����Q-�s�t�f+a4S��#9Xޖ�c�ՓӍ�0��\[�#p��PbT �5M�r��i��b��Kò� ,Kse<��8�mi0)��`VWDaY�a�e�Nx0�+Ý���]3�GM�a��\�XOh�|�Z.)��)�&	���$�+���^��E<G�^~��6t!�"� MR`5/�I^(�k��K��^�\�"T�����ޟ��-�yh�wv`��3�%��	���]�T�Y���;�7�J�B�<@��l�GpI4_�j@��t��J��縪dD��̫ ~��h�Ӌ��s�<2�V��o�":��JM�ԊJ�[�g?�E�6�1_ ��	�܈�[S�P���2��K\��5��6zcf���Η�c��9uɑkD��i]��z�Bm��|
>���=���' �J��M�:��'v��˧����G" -��]8|�<6�އ��38p�"v�M���@��_ٮ�����Q)�LHCfA1����WR������kx♧��Ԉ��|TVV"77a!����͛p��~�<y7n]��o���~��޸���ded�8�e5�+�@yI>ʊ��ΜQ'����w��ڂ��z��֡���eMHϩCRz�KQTс�-<��	�J�	iEH�.CXt
��rP�؉������y����i@��V<��۸��K蛞FU2����h�"|X�������U��F�Ȏ�q��a��C�}r?N�׾�86?���7���>��S�I�@�����>E��'��֓܏�/ɽk�ޮ :tl�GF�yH����� �yN+��EɶZT�[��;���[�?w, ��'��l�.C<`�	noA :�P���L�x� ��h������D7�XЌsA|�3�9tEt�3""f��`[x�[� mwx��,�Z�6�����瀀 �2��/��¥�(7`_�'�	�|�$�71�G��BY��s�z�@l12�ꡆn�D��yD�7�M4�r܏��t������D�������\7��D8I��_��JD�/�@.�s<$�a��gA�ބI���8_F{#(�!�,`&�#��d:����� �$#81A,��  �_E���c�����
��7�Ct�
�|x��#H��P����/��|�����5��e]?���u������P�{qy�c�>��}���M�y�z�����?�`эpt��������}�XB�/��r���E�i��$�D�'��MP�%�=��/%^I�&�{ʐ���������e���.|�{
�����t$�S�.S�x�S"A����������5�W�����-���%�N)|+qL�Tq�c]�'>�Ԩ�I�*#)I�J����ฅ9Å��S�-\�O� ���5��1�[�1�cc�s6�o���an�
7�N��>��ߊ���pnN�ö�hh�DL�=�S-��C��8�>�v9��eP�\��v������C!�������N�f"*�^|�S�/��Ց
��88���+�9�s����-y<GdD۪�pSXX	�0���.�og]�X�����Ÿb�1���Bww�c�,�	n��@��9��Bn�� [d�q�1_�`�5��F��R���}+��Q*���>0��V<���?Ț��F$�uz�?�	�2¯�?��ٱhΎAsFZ��В��$��b<Q��:R ��X74&x����>\�-)�°)�fWI�+�0֐��m.D{y*�s��T�ơ,+
�i��OEnBr�C��D3*���tC�'!J��� 4�ahx���������)�fr���h7FAK�ٮ��+�׆°,�W��?� ���7Tܭ�w��6��NW���$`�r*]5�]�!k����9�Ǉ��??ů�}�N�s>, j��@os.ܜ�U��X7�-N�fcuCB7�c��Kx�[o��＋7��|�w��܋��ѕ�"~���8��gq�����K�q��g��/��^ǫ���8������?��p��� ���'r�7_�j=WI��%5�1M�◠�>�I�of+�� ���bs��j/��@�'�E����ED���]x�GMp�k��j ��WA�@-���`�9�v�g�Ptӧ����LX�� ���~��w�b�#�>�	�;�ἣ	6s�v�Xߕ��):-IX[�5��XQ�u��0 ��k���2++���:�r`��f��`��f��Xח�u�0h"�saڜ
���O�r�Z����@���R�q�MEX?���t�OV!m['��vý� k�#����V� ��L�N�ylv<{���}w.���O�O��3_O|�5�|�i\|�a̜؁ڱfd��#�)�-�("B7��Ɠ����'.�gSB��U� ��xXG�4��.!���2]��ܰ�d$ug!���X���F�^�Ķ'vW�h??���=(;Ј���D��J�Hs�W�hXy,VY�Ã:�	ʵ��h��e�.��H�OG|S�"����(��؅.����l��
:�)����*=��3D�[��/�w
÷�1xs��WG�qy1tyc�'1zmӏ�`��ݘ{f6�!B�m��e���z��dy��<_O��\��j�K�HͧԒs|��&>v
S7gp��8��)U�ژ�T��n�̾}�s�4N^���]FC��R�Y��Z�$������2�M��3�۽u-��P-6�n���AX���46�#''��,3z{������HODcSه[��¹�簉8ݱ}���@Ok������L���`�=��_��?�4:;���(b���E�MHˮEYu
�:�rĥ� 4*�V�G�,I�)��-���ڏ��Ld�V!����QMlGs�����G�������hGA[b˳Yn��GJ8<�a�js�2X� �T���_g?���ޞx�n~�I���2FonV��J�w�t.���9�_h/:tu�ߣ\ӻX���枝=�����8��~U�������ъ�Yb}[���P�W���� mbY��`���k@�O�� t�šh�Bm�/*ҽP��z"'��DgJ�#��e��0[D���h�`_3x� ��A�,�@��i
OƔC[��!�g�Ü�B�3
��$Q�Lͅ�]�.D��ADW �%��@TrB��\�\��B-��� �Ǧ�&�b�5(��9�AF셱�����e�T
$��^��
cH	2Y/:)Q�b$ב��q���}	O
$������-�|?R3�������ss��-q��t!��e�9ȅ�]�1���nP���I
A8w�P�e���<<-�)��'}���RCԼ@��t(�Bz��L@�Gd
8��A�� "��d|X���0 #AY|Lv83C� /BP���徜�H$f0���Ov����D�k2�H���Fg���q ��́�'��D�І�t"d�=o��lKb�2�vġ]�/��=a��T>!i�i�$wX%��<��I��H��qe��+)�0�|���܊�C�'(���iġܦ�,�ˤ��[u��HXD��J:'
gB�#&XZ���V�&�1��N�6�־zp0�K�)��,��"��q�O�`OF�S0җ��6��>�%<.����@�s��O�M�\7X�v�k
�����|�9։;<�]>ӯ��&���r�}1�mS|{2���|_���a��8tb
c�eh��E!E�^�������j _G=����u�Z�0#T�b�9ۻK��?�,t�ƻ�&����
���(�C��ҽ��d��u�7]����C��)b���?$q��vBH��#�5�9|,ᄂ�H��8�OEEf4��ƜX��ţ� ��td���f �PK�V�x�"����Dm����tŠ�.�-m/� ��Q��ƒd��*B��0���(M#@S#Q������dƅ"%*�a~�"4���g�"<9�Bp�;¼��s�sZ �s�[�5�aX��U�qX�BP�m�R��>����y���w�������[>8����x�JĲa�7As�X"�O�a�X2hG��&x�2��Kx�W`����++�S��<���۲�|&n����Й̃��
$�G��8�p�k�`���Qvf�&�aԚ��mM(=�Cw���[����7~���������s���?�[��&�^���]]�+��4�+ź��X��D�B�e��Tj@�%��w_'�)�7�h��t�3"���,���,6qU\��(��<�� ����/<�D�D�{�c������2���^|��_�Y�� T�rh����j�-�P-L	P�5H'@�O�c��,~��\�����|���@�[�߽���w�=.>y�.BՑi����L\6V#�8)9��G7���NL>z#7O� xSw�b�����c/�6r�4��!XØӟ.��J���b(fq�������[����D�*��x!L�V ՛)�P�b��ꚎD�η�̷^���������<��L���IUƞ8�����>����ӿ�3~�������3�����?�/|�����%^y���-�MH�OE~[.��p��sx셛���l�=�Ȋd4.��*��YQ8�ð���:�[E�Z�ђ���\�NW�f��;�w�Ql��U��܀hš&����d�6T��Jܲ�F�W�)�.�]��y?@5=�~	@��Ȅ 57�4�5_w�>@[�R������Ǝ;�sl�K �A�� �G�a���\�x-��xv�·��k@�N���h7P� t� �&��J��a�_"b/`�@��E���7`��y�{��ًѫ��~��hz�x�[sp(5��l�>�S�Ϊ���@���������9��o^B��1���������;�K�=J|����nt�N#�����,u��t�MjK��q��i<��Sع/���Q^[�Z�����Ũ�*EuM9RR���c#P����H�/}Y�CCK=G�=F��o�ܼv�ʹ
˵a���,Giq1���ko��#�c��ndf#>)i�%L�[QY7��!4��#.�A�O���r��f��k?����й[$L�r�PXҌ�rbkhSs1��(��?���QTt�!���y�pI�+���r���9�̵ս?W�ha����K8���z�n��i<���ㅃ�<�>��E~O
�Ⅱ��IGC�������:R[� ��I-��� ���ڏ���p�j��ﱽ�}�������P���<&��l;�o�����Y�H��6l��І�=<;�ej�1R�*���=%��.	Ck~ j3�P�� Z�x.��BwZ�#�X���d�d�&���b���~"B����e
_�4(��Ѯ��,�δ�!��%�H�L7BJ��j�����D�4���y��_$EXJM ǥɭ[�<�4)%䈱�h���h��z����&�|~"O^�U����Ýȕ�v��}Q��H_{�����na�f(�s��v+n�q1��3aq_�\L`�b����a�h C�T�8@��p��BW:U⸑�)L�z&.�jh�ako;��:���K�� W8q{8p���;�&�Ŀ���!� {8�9s���^��.����
��HO���o�G̝b����(�����w�n[�z���uUC��\o�Y,�nir_�>�r���#�Uї@��;B?�z��8r��nt���-f]�&���0`d�����u8_+ё?��Xwo��{��/���>��m��G�2Z�r�QC,�d�@��������LӀm1�-[K3333333[l�d���b�)�'���p�'3��d`�����Z�Ȳ��9����}g�s���������T	��O5�9Pw��T�l��8h`��:EU���l��h��KN���n��xSDě!(ʐ>ߚp
ւ}���a�d
�$z/����>9�Ѝ6�I�1\�-�b���H�_Q�Ǉp�H?�$@�a7��0#���D��,�ٞ��E�@!��K�Ҕ�z*$�ѹ"7�Ʉ�@B���.������q�ς���m�
�*1�  ��IDAT*�AOA������ +d��'���>ci㨇({=Y΅��:<T�j�g#Uxr?QC���(�`�D?
�BB�f�@+���@'D��#9�ى�(LCUfsИ�ּ$���c�*���)%X%����Y���dtW���>ݵh�IGMm:*�SPX��� $�x")��ٌhd�"76�q�ȎEZLR�	���A��+�|����w;Q�'�u���3��\���Xw�$�A=�򅞐.��d�?�k�X��p��{�Pj�x�}����G���6�Vu�<�����w�A��J��p%����pȷ�A�)��^��{�9���Lh6�C�+

������h)=LN���ThQ�ca��ygW"vWL{��������A{A�d�cI*O���kG���!\މ���1xi��zKnA��A�&`6�~.�ytPe�ty�05�<�M�� 5�妴3��<��Sm�������k=�ZG¡ D�<=3a�#�ozܜ�����xd\q-��x��?�!�����_����� :=�4�6�QZ���� ]W�Y��jV-�!b;��P�vb�@��t�_e*�#����t���#~S���Ͽa���Xxt������uI����o�1~ģ������ߟ�k�������o�����׿��K_?F�p-T�B�ٞ*4�U���E[�~t���������CT��w�7���=��܅��^�ա4�j�=Rl�S_Ĭiŕ_=��t���1n|���e��4�aV86�>���-���k������>n�qO>�~�9>��S|����쫏�շ���_}�O�z���_��vc��*,�4�����r;�^>��׎c��OV(�R}aN`����~��2}�r\�� ���F �5�y�-F�R4ln��� DU�[P��9�ʐ��X�*n�˵��7�^��e5B���4d4d�>�� ��bQz1@yt\��EUC�Z��֝��<^�
lx��DT'��$�U1hߺ KN���*��[�T�F�3Հ�ZE�o	�QѨ�b����x�
�B�xA�����
��
Mp	";D �C ��!�Z����U76`��;6�Ɲ�h�Ӌ���B�'�nW��͑�+���f,zyzN�5�b����<ԏ������z,<�
i�w�GB�G{q��8r�%�,DmG?��k�쒊��l�Z9��PZو�����y���)!$�#%3	1���#d��#+;�A>pv&3�Z����i�(�%��'!4, �1���}`��c*x����fB~^rs��y�|���������!!9��NȢ�̣�&4���5M��
D%䣥k!.��n�����Q^ތ��|�,X��+��kp%6�<��/�Ħ�GP?8���zė�#(7N�
��r���\�)�&% �;-��#|�ŒK���N���v?<�����F&O�"՘G9��m�����z�wy�O�(��G�m:�Q�s� m>@�g�����a��ͭX�w �N�D}�y"���o+V7�pi2F	������\��xM5-+Q���I)%��M�ZN -_[)4� �[$ �!b�6�{�>�uin�HrBa��	�6H��B͑@��X*�G�"�Ka���A4��OՅׄ<�m���Z;-XN-��9�Q���#Z�O�Щ#���sa�
�	�pMDg����s?Nk=������K8G�℠�e2W�V��HSi�ãЪ�	#��ȴ�M�vZD#ت�
���6m�̣EYK	��DQҢ���g�H��V����u����,����Ӣ�<cdi�+�A�H�%����φ
�D��s�f6�5ZW!�*��C�TM���Ԭ?�>�ST-gC�zf�j	�f;�`E�^*%M�к��6T�D�Y����u�y��6�X�T$tM����y?}(�<� (B9؈i�0ƞ� �L}�fO#aY�L�)��M E��0����bh*�>
�S��)d#M!C��-e�6�#>�A*� ����׃��>d���(�9O��>n��%D��$d.�fA�QJ�jPp�Ϝ��<轰��\y�z8���c
�0}��ρC�S�`�m���\�)�:?�F\J1�uB�e�\��������	:���*ԀF�[���d�ü<6U�(
�e���{��;ct"j��DY~ 2��a�� :�{!���N���ׅ�-G���6T���6J	�=���04���:�y��Tc���!�����!�tn�s���Yp3T��|��R���_[#2����hgD�q}|l��m_;���"����D?X�(HBKMz[�1�U��U���>�Zڅe�ڱxa+FG�08�@?*�hl+DYu�K���?:Wz�;�'� I�B���p���(?dB��c��b���4�h4���� ?������pq������e� ;�1�3��N��l�;$K<!Q��ZH�
Mp՚����� (g��~���!~�p��{h]��d(V�S��u�C��)�C��P�Z_�^:Vwd�����(q�LC ���<�s�B���!� :� ��$(,L��쌀�H*{i��@Hj�GR��<<���`
4za<��|��e��3I0�I�yo��Ra:��9}�>g�e@���SRL(ϋ�Ӱ�����I|�h2Ԟ /@п���\)4�e�2�&�953��E��5o��%��҄H.���+��HS���(���)�*@�	��1{��K�����}��L���9S�BN��o���?���� =��E,;�9t.�i+@�*��^�3��G�����xB���7��%���|�o�a���?�����w�{t3��`Д��ḽ��MC*��9�/��<��C<��C��q�7¯���������"�L��h��
��*� ~e�}�:>�����_��G�P8�� G��a㵓x���.���*N_������܍�8��%�t�e�}�%��v^=��o����^������gw�苻���2�ف]7���t���w�?/���0��v�'t������p+̎���:���2���H_����R�,�@#����$@[�W�����\S�4ѴHZ����/�j@%�� �U����_tTG_�ڳ�9�A��GXe<�K#^�����	n3�RN�Ө�� m�B��J� ���1i{���Qh~[�S\lkAO�B ��jh!����ZJǫP��N�b��R� �����<7�м� �q?�ᗖa9au�˫���F�	�l ��ܢ��i�Ϭ��5hڼ ���0	�GHN7,����Q�څ̢J$� 65q���j����Z��ǟ��ɓ��@z^�ޖ��4�I�M�FFf
������	W�%��; *�����(AZZ�Z�����y�:pvu���7������!!����@uM���:�Zj����H�F#8"�����N�u/GEm2r�(�����ز	�,�@EQE3ҲK���Jl�{|�=��~��w`����؄��F�T�"0/�����y��=,�k��Y�		9	h[��Юe8��%,�<��7&0��.�ye�'�e���8������v�ܟS��B���#��C�	.�������V�(���:0tpkήF�0Q� P��Yߊ���H�F��A��Qp)�Pq��Mp9�ꍵ�&�P�������R]P�섲D{�� ?�
��VPK���bBo�"}�c�po¨B��i w=�����a>����bJ��5P�\}9�5V�\S̢���Rs��`D��W���N��� e]E��ӗ��ۦG� �L���<:�Ln�uy-y(�z�:jP��Bq�*�T�m*��O�S�Q��jۦGt;:i	��&�������U��ʓ��F���҇L� +��}���^9����S����Y�N��l�<ő%�rl�y&��s m�u�[͂�5����)�̆�%m�m�.G���4)sDK{Z:́��\�8΁S�e�\S:�"@ɸ3�Z�.Z�z6=x�Sd`2�3F��ނ~�E:H2��p#���	��4E*��HF�D�adNŦ�R�����Qx)I�O�D�|:�	3�D(%� c�@=¨��~���с��6d��zɸ��B����R9F)-�����B�C�޺С�m��l��Ԃ9�6��	ְ�5�C�� K�T��A?��i\}���5��O�t[��Z ��NĶ��ނ=�0� 	����1j@-*�aU�_�g�ÿ���ظwå�,AI�7
Rܑㄔp��Z��J�F�r�/���.�g��D���BMh}FZ2�P����;d��#�͈�X������f�h��B�PXj�����W��-�g] <]t��f� /D���������� �Z����^�p�0����c<��،Pd�$ �$��L�e!9��Q�4_�$��-�Y��/��u��}.s�tx���1�wFp��"<퇼��$!7+�Iሊ�%,�#0��n.�cg/k8�;�9ޛ�}}��)G�#U�N �$A�k@�j�B Ui��\}d�j�ިߵw�z�|rw>|��a��*��m
�Lg�0�T�"���HHFC~(JC��H�o�L4�)��Q�����T|�j@�F!CU$��.L�� �C�K�@z�pJ��8�t)"D*󈜉P���&k��"-�(�DXU_��Y�r|�T*˳����\���P^��ϟ�)��n����B��IHN�дu�ʹ�P�I���y�"7q�0:��_A��Jz�t����8���S��N��T� �B Ue����Ḅ���T��Ռ*7��ć�}��(@������#�cO���?��C��bp�Z$uT#m��?������y�������+ￅ�_|��_�������ۯ�凯�����ҝk���u\�{�>�����!jy3t��Wߎly�^���߽��O����^��'(\� �!Po��^&�5z#9�ݝ��Xh�#um'�}�:���'x��'�~�j��a^��*R���Y���Ǹ��..��x��[�v����c���;��w�"���E�.N,ġ�Gq�����.�~'�ƁS[�}��<����~����!'fy"��yN;�S �;���sa0��bӚ����	5�M[�0tjM�{Q��]h��?^)Ԃf�-���D�	MY����y(]� ߼a\��I����h�}<�����L�U��)4�Մ�����
38�:���W%@#��ro���2���XOߏ���n��xPn��}@��Z���[[�>�3�5;pp�?h��	���p�(<
n�n���`v� 妷c�Wa��
a���P��4�����0�.�Bߩ��9���a���($Uech�24u/@\F.|Bc�����4t#:>-�8z�4-Y���8$g�����ތ��l$�&"-=�apww���+�x�2'x;8 ;9	+�,�����o���W�c` 3K+�������N�HH�GhX����?�?��ϸ��ct�#(<~�q�LAd|��-����ʯ',7��y �c�PXތ���&�!.%�^�p�Bc�6�:�α�[�#�'P;6�Ȋlx�D�15V�>��t���=���N.�U����R*Sq����}�_�����>7���߸��<�^B�3���h:�'@�!:uP���5<[� �iXx"h���iF���ކ�]>4�5�֠s}�6�백���v䎉F��>���J�>���U�/�Z�
(7��ӰpP����e���ɠ6�	�v(��A	E h�%�#͑f��ps$Bc��`�h�(%���~T8�5B��!�>nzT ԁ��6�l�0��9WW:2P7���1�0����@͈g@�$�*��	��J|�Q�%tN�����g�j4	��P�#�Qu	Z:��&tM��6��h%��2�^�nO���������g
ߟ4Uj2�R��WVִ&	�3E���eDρ��K9¨�)�L��G�|.�$�K9�'�+dlgCƎb�),�m�q�R��V��h)K��mv� �@�98	��n�4%��B�IwmHzh��i)�EȚo�H��A�0&��li\k�l��9t0]&|Jv	y�@�(Q�'��G��� � X>�R�O�I��؜��ih��� �)�a�cH
�uF(�Y\#*�G�׆P)�N�v��FK��ȸ�6~�]�A��H��2�S�� ��fТ�>��@/��V�M �d8��Pi�aMp�!�=��0�B�'Bd�f�L{��u]	�1Q��[����!.���W�����Z�Ü�iA�
,D~g:z�֠�-���h��ECi
R���(/s�����	|]���hw{}�9�����PoM���ҹ��q�(��� k�c���ڈr�E�����.ƈ#4&zY!����pG�iÏ��sփ���Q���11~V�w5�?����^p���Η^����t=��Т�A��󼍡�g�yf��~�6Љ��^��0G�y�/t�ܠ_�����x�:�inpKr�G,f� {�:".6�IH"|��""� �	�@�	�t��$���k�H�B"����*5���5�e�*օ��@�T@9���:p�����5��ޫڱfY�P���B{�P�)�)<$�K�d��r(2ñ�%TJ,���<�Sj�k;����;e�"E� (3F ]�@ L$�18����Fy}I2�.��5��ƒL�,�yZ��d(�$�y��@Rbq��4�,˂ʊl(�y+�N���}3g (�k3���iJ����B��7M��PF(݆��28�f&�(�K��D���S�:�Ut!�à�	���l��# ��M����@�7�B�6	�YPm���b�q\*`�,k��O��@�����N�m�r:�ѻc�|�9��_���op��8x���־t�/����	߄�'7c��C���&���m�yr���)�����>=Ӛ�I�AԂJ�{	�}���x�	��޺�sｆ�ﾊ��[�9��0�φ�p.��S0�9�J����/}~��}�>nܻ���ݘh��4�}�"�&�ޢ�g��{eK�07�Z��0��A�3�5L�a���*y�,��}	{.�Ŏ[���z�޿�`��/��kdY<4�Σ���^�/�R�	��O�V&L�Ӓ���l��`q	���c���蓼v7*��Z�\���&�k��~�iKP��	�t�ԑ����ՠF U!�2H�	����H�Q�� 54��bcQ�<�HW�G#�:�%���v�P	�ƻ�4	�jB�P�'��vTmj}Z*������ �"�V�h@þ6��mEŶz�m�C�D=*��4;�H m�4�%�����@)�ܓ�=9*���|��J��;ԍZz/��a������՜	�xO�'����׬�����,�@ZN*k	4M�(,������?��Wa��c�N``l=}�m�CZv:�2Ӑ_����@X[[���	�.�����B�}�Z߈�}ؽw/�O�a`l
{'7�Z}�����D��
Ӻ|���8���HNυHb�r��^L)ABZ)A�	��HϭCzN
��QQ�K����w`�R�Y�и$d!!����Z�
�+� ���Ip�
�U�7�Ǹ�4�F���4��;�S^���X�k�=��E&���.���݇Ѳ���޴(�����y���)�*Ԁ�J�q����FB-��D�v�l����!����!bt6o�y�4u0��!��\��|h��
!��*P2�(�ը\_����TO���t� }:h���QG����Ԍ j��s$B�B�#6�
y��M�
 ��#�>B���;�>F��2�|=L��j�y�7U��|%h�W���2�	�\�uCU(ҺaTe����2]�@۞7I��
����(B��)��$,�XJ�\[�
y}>�&�V
�Gy]�R�J0�m
t�h;m`:si��~���*|���t�L)��$#��e	�S"KQd`N�<׌2B�D�u)]HͧcQ�L踦�J��9��"I��:i���H�4m5�H2@�@�A�.�v:�r:T)R.���<!��� 15SB��&*@s|
�	��P���HЂ��S��!x�긶S&��S"E�cxN�G�kB'#-������_(E�����Is�k�!��K �*(�O)��ȸT��Aڙ�%O}�xB�@��iL ��V�%�=��B�G�;�;�]�<aW��g�O4�m�#l��a�b��)�0%|���2l�NKhMG,�lm$�6bצZ�I��p���e~�/,�DӰX�x�#�	T�I�GB�+r�=PJ���P�d�!9�an�p7ׄ���	�����r�owca�2;s5ؙ(!�qR���N(�rAy�
�)^��q�G����D�%!�kA����VH�!��Rm�d�X?KD�й����o�x_k��%�=,�e�@;�;#,�>��0������b^�54C�� �
���#2F�@#�j�vPK��F�3�f{`N�ԪܠY�yU��#���k_��\��K��K��	�~�p�u�o��B��솀O���+�vb��=�>I��-
��4
} K�d���I ��˲P�j?��B�&L�*[ٚ H$�"sE#nu�����.���`~�k���DB�'\4(Eh�;� �ʣ�J�R��ܖ�)C0����kJ�c�0H %8�.I��TH�&Bra"�&���<_%������JF#!��)-K�
aO���@��#���R��+�$�fC�P��'�	�< ��2Q&#Lhº�QK�2��S�
�5�eT���
t���B	n\J��	t��আ 7=��0�Ġ�uyB���~u� G)z�Pq�ܩ��O��M��s��8ő��3=61@�y��g�9=P�T� �A��/���Bm�AɶnT,i$]
P^N�t|r�cn:��;�f��5���M{�����w�;|�C�r����	���w���O�淟�ܣ�1vl������)p�ΆKW6��P2� ��_µ����wq��������o r���K.��*������>�������Wp哷��o�ĉ/���=sJ��K��ȅq_:S1�4q+[p����������'x��T-�¬ xT�`������/���Oq��w0vt3��b!`J�B:&�C�ʊ�YI�P��&����>Mkz���&�~���ġ�q��&*��Ǣ����g��� ƄP�<̡��PhFۂ�a�A�|)��H���-YVN�v����Z����
�e�����+����ʅ�q�W"}Y*�6ÿ� �+�� PU����d\���� 5�o���0�с;A"�<Q5I�-
EHU�F��<AP��������@��4�L �~�P�+�v�ߧ�(���L�>��PF���F�h՞�3>)��^��	e[�QB-�҈��#��p8���!����qy$\h�!�<Hݑ4�@�a�͉a�� ��^��kQ?���(�D�"03
��V��bl�zW5������B\|�:~���� :g����M
RTZ���!dd� ������3"���i�ù:psp��|3��օ��!,m���/�@89y�? ��񈈊Ƃ�!��Ʊ���%L���M0fpV!2>�y����f���Z�4����=�<�ቨn���7���{O�~�>��X��%�Q1Ћ��:�Uf��0�YA��
�x;`��T�� E��$�45����XvnV�؅u��Ų+kѴ���zж��:�&�S�)(#�G��S��iP������ PQh���(�۴��7��gw�_��q�l@۶-@�dP�k@�G�iX�W�� ���NN����)��4,����B?P��!���E[�7�-�^�NrFE�JblQe�J^�r"-�MɊ�@%��b��`$�!�NL�TH��#�>c|��e�}*Rh{X�)��M��sK5�(Cg�
4����M#�)!I՘NOeB(CT�P��Y}^�B��&��G�����DƦ�ddi�E^W
�!�����j@�k;��k;	�S#l�͟Yz=����rL(�ts�賑�"�ZӺ�Ԗ�jǵ��HQ$����\���#9����)�Mk)�����$8�&#�;�T�N!�#H�$'#)^�u^���,e�:�l�|��d#M C�����|�%�h)cN$�NOt�HǚC&�BX�eɘ��Q3�!̵���d����*I�
������k���2u��"�K��(C����J<p��T}��k5�
" ��B,0;��>�P�цU�B��T�o8y�6ߍ���G��:�(���Vp(��[�5<S�P��uع���$16��DB�G�� Y�RO�����2N��p��F`�R��J�s_/c$�;�,% 唌0':X��v�����Q��zp�2������Bu�sSe8��0��Ɂvȉ І�"��Ѯ&w0@���-�l1�6z�r0B,4��N�Bhr�=�'݆0�c)$��ᾖ��']���EP����	�_�E�A���D*9�z���N*�g�8�ҝ����,�f�@&Ǖ��|�.��Ny �˃aP��`��ü8�A���uN �R}`���D8���1�t޵I��5�s��QF��:F���A2���ΐ"|J�yB��K�Jo¦jE}@�JMI�|��v�ɏ�O�->����i�+4�JMA����h$d&#�Mp)�M�/B�fX�����*9�Wr$�#�Ԥ����BN�3��ZJ)�#�5v<�##Q���.s��A'��k'#��$�>���&�	�%_�A��?Ef9C�������" ���Qd��Ar5=��9�$��cPƵ���x*�󠲆���\h�p�U\�� %p�s%�I�!`ӱ�h�����Jz]VF9�.I���H�k!AǑ"@J�c�&DJ1@��"�؝!�
�@��_�Y�o�W��/o�¦��b���B}S)4&J1{c�7�"`{3J��rU;v��O����0�_'����K��Х��5�kfD)�6C�����r:&��������>O/����%]Ż�s���~���;нx��������<y������W�"sM�{�ຸ
�2`2����0hM��P�7����:�zp���%>��q���"qI+����W�������}�[�<�+�����7q����g���[7	/c��V��n��ˠו�9e�ZԈ�t�����#���!:�W@;�v	�x���<��K����۾�b��W	m:O��9N!�JE��UF��r�$�t�W��׎��s8va7����[q��n,Y;���88g��8:Y����
�TW̎��V�=�n@#�[N��9ك�(Z\J��*�moG7�����h7�v7�t[��	-���B~�֔!kurVT���+a 		(jHCUC�@�@ UƬ��P�P���
���:�Q�:�YU�r��l��h��P�fz0p�߸`kg �4!Ea���C��:�n���4l�AA�l}OƛP���
�u(X[+�׋�s�-!t#���:�lt&�PM�!lr_R׀
���A�6\	�\ʰ�׀%�L�Z3��������N��R#�n�^I �yU��0D	-{��z�g#�QC�y�Inz�L m�m���!�L8�86���0rv%���KϭG�X%R=��k����/����k�0�s3`dc{7����w ��~�������k{�G���
�׮Dvnl�,�lmo{G�x�������`�o;[*�Y���	n�p�8�x���>~HHMAlr��ك'�~��[���['w�$�#����Y����)�DXl
��j�YP���LUu��{O���6�j�P�ҍe[��S����{t.<��5���V���x�F�)36�~0K��I�t�-�i�I	��S@qw�\߇�w`��8v=>�ß����KP�����d�pI�0�m7�o�~����`z�趼�~�-�lz�h��Z�m�6�oC��M�ZP����؀Ν�S��A��7��h=�nG-XZ���"d�#w�sU5A���Q��R��(���iI�Gn��}A+x*�-�T���� �s��L4�{�*�eq(��EA$�NX�P�g&�3�� M�"�Z!%�j�DS$0B�`�m�h$�3�
�a��P#�v��� �n���/����j`!s��� Q5%�(C���q�P5(�(�u�&��J�N�S�NT@�$>őץ�g��ψ<��{>r�P9��26g�t�
�O *c9�VkM�2@� �9�:�ՐN"�#M ����
Q�o�� J��0>%x�k'k<�f4�G�NN@(_7-\�(�p�Ĩ�"��C� *K��aTN��d��#G ����r:B�gf��@M 9���;=^���	�2BM(�N^�O��'��P��"�v
�Se}h#�ZC5��f�b�y���fywM��σc�;����]@�w!6y.0϶�q�%3�`�K -��K��2��2���t":J'���lI�J�����rO�T>k�h��:����
~)��)�E	&x:�� [��x� �ɡ��q҃5}Ƭ�VNڰ�s���<�aM�]�Y΂��*l�4�I`t5B��b���a���w6F��Blub-J��!��(�t2Fa4�e>]��6A���6G���,`�e
np�'�"�P�4�=T�rI��J��B�#R(iNP x�e<�݄>��V2�
X��� *OQ)�] �k�a\��50��qE(L�"`Y	+Z�(�%-mk"a[��p��E��%�����^�%W��J~K7H@%+} Y��o}	��� ��{-CK��PȔ�@6��K�p��U|�����l�cQ �б�ZC!G ���D_(�D �I �%Gf0F���2<��:׌r3݅�$lJ20�D���}3���Ƞ��7���Az\N��M2P�z1>����: �8�K(�O�eb�r�WQD %�	 e\2
��0@�	f��!C0�$�����YP$L*��Th?�5N����v����d��rl2ny��#�n����P���=z�x)��$�1*G�|>��@ϋ��#l��J U�H0��K��>9�K����7��k3���n�����~���51B���<� �|D��������g�?�<	��>�Z]��dD�����y�&�lGˢ~�|o��3�'���۸��=������nY,�V�rU%,���au�	[Fm��\ьMo���?|�K�~�߽�Б:�&y"x�
���ƽ�~.�%�C�~��C���1^�\~�6&��D�V:%¸3�����bVqB�jp��-<��+ܥ�v����_I ��un�^9���������w=[���H4��E@�`8�2
*eaP(	��T0��ymV��C,ݘ�so^ĵ7/�إ�8tb�݌'w`ņa�ץ�=�
�E�0$�je�C#�s��a@u*�we$���M����A�p>����w_�_^����.U��� � ��W#�
�Ykˑ���+��� I}iH͒��y�ϒǜ9��O5���BC]ʊ<�,�Ty�!��)/\f�r4h]�y�3��*�)�A�a��-���,?DTǢti-�w�u� ��Q���$@�g h��@�i��:.hՖB�@[`�kV����`�;�������#�����l�P�r� �J�+r���;�C�'�
 �G��atE��Q�Z����ѵ{I]Y��w�U�3<����Z�MGv`��C��ʁ�'���Q44�!/�M��(�,����C�V����R$�%����6p��E��;��6����2���3��[;'8�z�U@�\��Ԝ,:N��څ�>����p��op8n�~g/^CmS��{��
w_���2n~1h�X�3W�����3�+����p��%<��c�t#�W�r��*N�[F(��`���8O�8c�#�m5e���<����>�y��/�Ǫ��qớ8��Ut����U����e5���<�����0�mj��E<�Ó��6Ѳ��S�V����@ʃT��yw+�,XK���}�Xy~�v@	�PD�PH �-F֢h� �"w]
����R��´,�w���e�B��,o§�S�P9	�B*��S7/�
�@�D5�����B��J_@1Bg�.�(�Z�#���k×�{����E�z��ւ�|u��W�,B�������ƃ�D	Yʄ-EZ2<e�� 3�O%����ԂN����� ���� C���	1�L�1�'��@o���H��e��0@y!�4~
@g��M�����R�n/l�}%g!�!:%S�/)AT��*~N����j|�5��ׇ�C����B�5�(�@�W��QE�0K̉��z�!T4�7Ջ�%�@�{�Í`�j�BOX���\a��K�y�̲,a�kMP��K��2,�6���t�rb�vt`�X2�}���
o�6��pl��gS\���Ꭸ�p��h���݈�����6���P���8;����Y9���� �t>0��@SX���6�����P���4W�u8�i��� ~�Q�f�Q�LKB��ul��@k=�����V��t.q2������s>ܼM��g
� S�}9��#�p����DxfC7�Jt��I��D�$S�EIw�T%�	��."|r?�|7Qx�k')�nP-����`�Յð� Z	ӆh�Q��a���HՆa~]̚h{s,��`՞���W��E�P��j��0ߧB�/� ]��*��3�uA��>���'|J��D�aP��"!:�;�_9�{������c���8�����!'4�%�R�T\����5��|��Q���s,AT�9-8͐) #T��9 �3="|<)2�C�t��\s�5�0n.�:^u�2�OP�5yP�c�̈́�)Q ��1��eWB	|���x)�z��O��9|r�������\��ׂ2(��)0��)P׋��a��P�q(Eu
@�n.�ɖJ8Q�"�
*�{��p�����	��ZP1@�	tc|����7Y����o^
S$?�7���[֡b����o?��?��_>�_?A�޵�k΂�X�V��lm�/-�	�lVV�jy%�F�`� !K���K�������/�FĢF�|xw�	^}|���;���k��������x�ן��/�C��Q�&¤;���S���F���|����7��ڣ��X�p/X��`եc���g�G ���-����<���ZI4�c�^y:�(�avu4�i�ؖ\��{	7�_��+�q��69��Ol����&����2? &����l�0Lu�CQ�	�������\��pQ���W7��d��t�ZPNx*e���63�j���
��*���
e+P
%cE�@�դ��*��j���
UeE�VW��*�75��&�^����r�W����$$ �"	�9�P���<	(��C�MN��(�g�H�;Ѳc���fKx�� �@����v7��T���ePB��Z��'�4�u�T��\��5���e�r�h��6���<�j��.�$�^���t�G��ut}�c��J�R��#�#�A�T�G(}��[q������}������!�w����a	Qp�ALZ"�s�[V_O899���	.�6𲵇��9�4�a�kkK;��;�wp��������	;'W���".5A�x��U���޷ �su`�ꉃ�Oc۞C�-�DFn1���=�H�j�����M(��Eqm7*���6�ë6`����;��\�Ц�(�kD}_���PG�P���)�v��v��*��k�=Ͱ`�B�x�0�_ق�s����I\��:6����P��U�����"��+<�
#����@�ex��p��^|��҄�]�h��F�h��G���z���a#O��Mq�~�� ka)�y�+�N����dx�� �p�7V��c��Lp��pt���9��ůNtBU���Pk�*�q�91\�a��hkaTܬ(+��Y#�
��d�gR���1�nZT��?���<�������nw*t:Qa�֖>HF��k8Zzj���Um%�U4�L0F��D�S�NF�Щ�p��?��/h��$B	��F���41�8b�Ғq:5��A�B�Jޟ���M�jr�,#RhJ�l�8H)B���$\� �h	ia��'IǙ	#tZDǟ�)��%%�	�H�1BE��[~�Q~=&1*K����4�\J�Y�Ќ�Ǭ'a��8�O5��0'�B��z����b��Ϫ@xW��\��r:q;Jm��k�4Sx����;{�4��٥8��C��H-��3\`Q��*��� �;^Ua�*	�G�7����� az%g�_P�3\|�0�>S��:��C:��B;��A�ho��a>!��I���`d�CKu��j��ANtLwWC�|݌��6n&�7������I8ut6���1�}M`M���)�8p>���1��1��J�GX~$�+��X'��XC*���I8%�� �E��!xrs�\7��A�"S���H�@����^P,�<!U����B�2U��)�V�/�+���Q*��a^�/4�=����[�D��5����@*��I��٢��W�p+M�!W�Eh�&J�T���L�7dj�������l�خl��{���]���5,�5�|��gwD� �>Y�)��Oq��$<� :2�'ta!��(�P�(�D+��?�fq*d6�D�IX��&��2@_q�'�S����d��� �M�֖���S�#0�����P��.�h�Ti2�渓���Pn�;u���� ���ZO��,!Y�PnB;=/��%���K���9��M��� :!��1�v]Rw����rt���7o���"P�1��?�%�	%�����T�<���� Ó�W�S�
��\������\�Y���t�(���s����x��Oq�wѼg5�:�༨
cePh��U��_�T�p�UGA��@� �dO(�zA%����l�D��6lz�%B�g������*��{�����������R�'t��#��M�qC
�۳�����x���?��/?�+ｍ�mk����(��|L0��/>ǝ'����	�5B=�e�]��P(=��`hT�bnq0���I8��9���m�}�0N���On�ɓ۱j���a���lo>u�n�#���C�b�E�-�� ����$�>���޳�K/,G�q�@+*�.�xAn+�n��	��+���U+�ReCEH)K@Z��(�'7�UU���,dd�r��`�L�K��`�d� �� �*%�P��%C%�[و��;�CG��eg�����-��� ��n�F�x9A�%[��J�/��(C���L�㦶b|r�g-7�jF	>{�Q}���3�{�6@׉��?���W��o�\ߊΝ�H�N#����j���ׯ��[�c��]شu+��Z���d��#&=Q���)+@aE1���,��7Gx:8���)Q���M�����vv�Sg��{����n������ �ڑQ����\�~?������w���������Č<�=|
?�����l�6\��6�]���%ȯlCq]'Zc��q�۳k�o��U(]Єĺ'�� YapK�k�/lB�`�aFNQ����4A�����Q,��	�'�c��]���{x��+8>&@����0B�&���BM(E��c�و�s��R�㕎)ܖ޿:������
 ��,Ԁ���}��M=�^�& ��c)Z^��Ee�Y\& �`%�G�]]�<������2<+7֠j���Cea���EK�'���P���MrA)7Í�C���N
E��(����!/�0k;#>�	��I ���F8!4��Bh	t�*t��h��U�
��F����bo;k}��jA� ���uF��
T�JO��!U�P)�L}��� ��
���Q��d�.c�E �q�����2�|�9�cD��?�҄��a|�&YO"�J�}Rő��:%ӧ`e�N6�}Z:����B���p��P#�(��F�@*h�@#(C%����P��j�T�M�<���ch��@�^Ke�yЊ0�U�3���Ŕ"wxW����.��p�0�k�)�3,P����Jqlo/��[���\�g:�-�P�f+B�C�?<"����P8y�:�F�03�S��x�i7��9A����6�㤅ٴ��5��
�Z�W�>:P�х��.�x�A�ˀN�:Чώ��\��g̐ng�W��l��p�6����	��>&0�s����}��`-z=��'��`v�	�M�j�D'��R��$�5�p/��V�d���PgHD%)R���I��R�)�����}%�XA"����9q��!]k�Pz���%�R!f�����m	´�;}�=h�I�s!A�9	KH���r��!C�Q���\:҂>ö������PO5ד�ݯ=��I�y���Z;H��%b���d\�w����x���X�l���J��9=1��%�.�}Aŵ��T�ʙD�8S��2>%@'PEsmN�x���HȜ�|VџP��#�'�s����r�-7VX�� 9@ƿE�:��K���J�m��$`�00i9=�U�u�eyB�AqF�n`L�Aj��g�j@e	�r
�vtL��9	���sJd��(]'(�����T� �1Qí���X��	*�Y���c8}�0��7H�o��?�����{{N�	e�r�ə���o(oetN� P�'=G^�?��8{�2�#���.��Op��wp���(#�9��¦� �=�Yݎ��AM,���0r� w���	�Q�yr�!t�N��0�Mj07�9��?~�_~��߼��'�cp�Z�;{ W��ǻ_}����n��Oc.���a^�
ò�-n��7p�7� ���ܵzQް$�n�~
��|�)���cl�z.�i�H��,(7�U��RY�P�R-i������1<��.�9�Sw��b'�P��]���h��]����0��v��D�B�ʛ69��@Xm�[��ӟ�"ht�vvb����R!� Z{��*h�v���zl�Cަ�l�"�֠x��)^��K�$L��U��d�G	F�,!���4[�ʖ�m�}G]�D9#�&��0�s1֟݌w��컗q��U�x�$��;���������8�^�����҉�M�cBb��O}@���W��k8��O�(���r��$�r{3��S�'#T�e�L"����j@	���]�;D�b�����0zN/������+�o�ؙ5h[׍��X�G��*�v�NL
C~M1Z�ڱh%�u�"4��"9?S hJ^&rJ������@x{Q�� ���`Ol]�A��m�
KsXZ�
Mp�>~�BP+[ħ�a۞����ukq��w1�c;-FfA1��2�������4�ԅ��3����P��C�ى%���a�W�!����X�}�&6�u� �Z�]��вT����5#�	ް��c�]��'J�P����
��1��~���#��b쥵���8n���|p
�GQ����ͨ��*D@�$D��P�'��12��G2�%,�jB��c��nE�nz�	����N�ނh��^,9�=�����w��Van]�K~��Qpg�'��[��:9K-��;J'��� tP�-����4��;j�]QE��e�+*)�T�+$�rMhv�O5�B��I�&p?PJ��� �hO!��ڈ ��XB]��<A�Z"�R\t����N��78���JFF��U�,B�CTO�Je^2>	�J�^2@�tG�"'������'!*�?���z�?+3 T�l6�,�Sc�#�>Pi!�PMHR$&ã�J1@�΅�o��q'J���#=%b�J2D %hr�� �O�"`��+< 7�j'k3����\dt�O��dx���C���Mg�.3g
rz��6\�ə�S�(m�����)�xZ�<�!����Ӿ��s����&�~-d	�r�J���P'hF�A5�jQ6P�E-�B@�j�	4�͠F�Xe«��6T�1/�f�6p�q�ģ��yt�'|��[ 8�5=��X�;;�ok��!� �G�d����N��A��wy |�B�Z��?D6� �>1������G�7�����J�Tr�E�ِw���P��O%����>鲲�4�s�ᡍ9�z��ч�t��.�	�:�:�uֆ��\�`L���1���1t�C;p>���,B�=Uz��j��P�σl�)���t�r��GpI,b�2�U�h'(�9L*� I�4�;�<��v�}�HBf������$�	�tN�N��%���b�`h�8a��5T��`�
׬(�%�+?�	�pϊF��~�=����F��2,ڽ���@��n8�`��Ql�w�M�Р�ܦ4f����e��Z�9fE�	ʚ�v[�ѺY�R�p��<��>*oc� jE�w�Wh�DCq Z�'��4Ó�a��Rj0
RñBD<9��s�B��`|.I�$�PnjK��Ɯ�g��g�I,I�)���`C�.J4�|�Q�yf�Y!����F�p�L��0HP�py����<���\�%���i��M%� D�W������m�g(rm%K�k.	}�瓁��ˌO��S�CH����xR��'�k;�֓��4B-(��+��K�A��6އ��2<	��	�3�ʄNUz�j�ˡN������A� j��~�u(98��ck0�g���gɿP����7�(�L�T��o�L��)/��iߙ���ϊ���o!Z���?��o�����([Ђ��l�|B���������[�v��d!웳`\���E�8�����_�O��������{|�����~�g��u�S��ӷHY��$w�a���诿�����>~}�W¿,�K�p����p���8��e���Wc�+�`F������u�2^��1���׸���۶F���΋����q�W���|��N�]Q<�rC1�*�+��QI��rU(K�Q �Hk�&ybݩmx��G�J�3�����8v|� ڇ��$�D��&n�Q0����=u���sQ0�cJ��5%!w �#�(]\���Xtv�O��������ă񼠅�w�5��*$��!�9&���Ж@Xv(��،ơx�z�!�	��)����A,?�{o�å�_ƍ�o��g���{������a�y��?>��Ob���]؈��6>7b��R��^�����"tVl"�"K�� D�2���Nq�2�h�?�Z��|�1���t��-��D��܉z.�tc�0h�D#jv���H�h��������p�#��h^'�Z����$��TTʯ���Z�r���"���l���JD���k�x���'���p7�_/�x�Vz�G�wz	�Pyi-���	kΏcp�B�ե�2��A��p7$� �$��M� ��#>/qY)H+�FVQ.�b��@?_x:;����>�X40��7n�����-��Mo�����7!��?)����c7�����׿"P�EIm��RQPY��z�{h�z	o}�	��؏���(�i#(�:�k�J����{�2���E犅��FTE
����0xd� j� o���s}���#�9+_ڂU�v`�K���V�|Ʊ'������Z�J�g��Fz��ۛ�VL6�ׂ����3�fG���d�j!�nw!��`J��$ ���2@��^��ݣh�܇���[׎�5�(XR���"d��<m�[��R (�����f�x��}
��T��F��Z*O��c�8}y~���FG��R=�£�fqͨӽ������.(�w���P(3�a6B-�0�$>9���) ��e$(�ݴ�2!�PZ�R3� L�� �yt҆��>a�D�>���n�����Cc��U����u��� }u��AEGQqM��.�"�a�
��wT��vB#��`Hw#����Py�9����T����OzϤ�M�"M �O!b|N��J�q3SƧ�٩0l�$@�_� �`�N�mj�	sC�VHqJ�I��L�9-2I֐N!��ad
؜���?݇kF'��F�"��?J����82�p��	Q��P��$LYC#����7'��h]����a�eui�|��|(�|���]:��!ۙ�腠� ���!���̬�@LL�b��V��X�Ջ�PW��� d6�!�#�]���JFvg2r3�7����l����Q9Z�����x@�V�\�I�s� ��B-��o�Y�yP#h�"d΢����o]���D����3���!f{�H0��:?]��h]��9��l
MB��03̢�s�jv�Hs�FQ�u�C�4Ip�c�/B�cW��`*L9e��*3fy�0)�uA,rB`����`Xe���~@�˓��]��M�X�o-j��v�0Z�/A��J��ބC�^�+=������7o���kx��#|����������|�nQa�7T�VO�-gy�?�:O�>�e��3|�o1qy7R:󐵠�˛ѳmC��>�а��{Q��~7u�o�Fv�`l�0vQ��3���e,=���P,r�Fw$��l	��Ё���,�� P��H�0ʭ$���L��DH,M"��>�Vhj;-BM��ʗ��Z�gk49b���9}��axN��MB�sa�>�f�B�XHy��(y�Q��"��#�*�T���f�|�
�8�'������t�F��* t������E}A���j:����Ϡ�@iQ�&�Kǔ^� ���v���2Y�����f�D	�je"���
h@��K�A�����T�]��{�������D34���W�?�Ɛצ�S�r�e��������o�}g
<4������v��M��}�!��ي��
��Wa��3x�7_�_|�������A�����.�Y}*4�揟����������_��y�/�w?���?�ۿ�o��+*�C'��t>�u�
��k<�����Z6-�mn��k��ѫx� y����u׿x��ｆ��J��F"kY��^��1���t^z��e�`� ��X,��7�:�3�����68�&B� ��0�*�S Z�B?�DYC'�	��������;�p��^�6>�� ڋ������ʞ.�a�"��@S�0��R���h�t�QH��E�(-@ώ.����'��(�l�mcrה�����(�҄����-E�H)�Gʱ�p��?>ĵ�_Ņ����G7��Wo�֗oҶWp��i#\�[o�ªK1vvO-C���=�X ���e94F����D��Q��B#�n3a�J�,��HH$L>y�[@�� ��OP��)\�i�|C� Q�'�	ZM -YO�sS#*6	��G���� z�k#�f��ȵ�{y�[�0sG���h��ф9���)`s/�pS�x��!`��˦�\�I�����#�hf�RxJ��Sc|i��˯m���m�xuzv"�66ю�	w�'}�#rb�R�����V!23	�qH�NC~Y!�S�?/Ozy!):Q�!���|��������ps�����P���X�y�e�F�p|�Vo� ��=0K�n��Sg�>0�����ـM�b��3�q��"���cK�t�vmX���Nt�"��IM)M���+;����N��U��=�\f��Y�3�GBC6_߇�7v���b,�����Gǰ�m�y�׼�;'�9-B����NG'gz��PJ���y�����A��3Ѹ�Yh�˃u�^���Mp�&z�0�- �jmT4
.B���E�k�U"��-�x���R%��k?��jPK�����2:�,*�pa r}ћ��L_��J�ѓ��l��{�� Z�䊊xG�#�� +� J�ZPn�+���r�g����0Byᦇ0Bg(a3����a���!NZv�?{�;2B�G�rև���t`b�=%h��ACK�O5B���
T	��t��H#���@_йB���B����|r\����)C����� *��4<���Mp�(��q�SanLZ�`B�w�J6�G�c��Ƀ�+rq�d��F"f��FsZ�ΰ/TF ��3�
Ȝ�$K
]�8����N�kGy����K��5�+��R�#d��@=�JQ�*h��cV�h
u���c�Bj��fL%؄b�c̦�y.�^��nN�����aHl�Dd�򛣰f])����㣸px���cbs3�mkú�=�|d;��w���?8�m�h��j�Êm��NP+v�i�	%��	Bta�Z��ݔ����f�>�&��~�cl�3�?�?�f�)�����L1��s}��E�:����� �t�ya����6�t"�e�G�:	яu�G1Iq�E��R���H?r�H,IERY��s��\���Z䍵"��ك��^Շ�}���,>�	�l�ąT {����=>��7����o?��/?»�����G|Ků����o�ݏ��7��%>��״���������x�ѻx�'x���8q�4�^y	o�O�/��m��Go����k���=K���V\{pw޿�KwN����p��a��u��Շ�����<�C�w��+Gq퓛X~~��P+��Zg8dD@b�G�%pr�'Óօ�����N�S|r@�$>E �Z��a`2,�����������z��(�rN�@��tߌM%�-\C�$�	S�0i��(G���O�"Q�˄P�	�J���$@���9�O��5�B�&��_�"T�ੲ�Th�����;+1�jD۝ƫ��%��0xtVY���1q������&j~+(Í�0��O�O������#�?ˋ�f�w�0@��?�9�e�������νv}W ���m��F�|���/?��/���;Q41
��|X�g#re}�:��㷸��:?<�[ﾃ��<��ܸq�����o���W/�|��2B�Y��O��_��K�G��.��og1z�l��'o�̣������+z����
�:��ԁ��~�)|�)����6.�q���"���n��ջx���t޹C���Ĝ� ���P�
�geJ�\�G�ŶЌ�C��Q����Y�'����G��c��^�S�;�,��!p)�}q ���0?���p)�oi8��~�ZR�?����R�/.A�x���h:�t��PZ�w���E�y3a�yO��a��2׽������'\�{D���w�c��ǰ��n�{y�Gc��B��C��a�"\B��^:�h�Ħ���^��~���G�Vz���"����M���-� ڂ�M\�� ��Ѝ-�<�<'h%m+�P�J��榸��Z�z�^� �k>�	�x$�gk@�h��FT��S�-#�T�e�(��7�mel���}h!���Aۑ>t>9]'F�n�����+���l~m����/GRG&�`�O�Zx^�sc�w:!�ψ�$�#�0�i�H�����3B��������(8�����R7�u�w��}����A�
Ext�s�Q\U���V��~���w������X�z�����`���^��ǻ���|�5ƏE��*�иxC��h%x6�"�&�����
�{z(�2�����g��A�DEhv�堍��bl�y ��ǲ�Xven���O.`�k;�wpj�6��P��]3���N6í�3��Ԁ
�@y0���r}wx>Ѧ}�h�4�j��W�7֣g�Ь\���)J�0Q���,*G�R����)@�	�r�N��d|
YW��uUt�) ][��%a��p�?% �فX@�L/a�#����KpAu�#*��Qi�l:�p-(��;u*�� �~��^ƈ�4F��!�]	�.�B�9΄P�g(4�QK����A>!/B���Q�N�p��;����2t�e�6O*e-%(k+C�@�B����#�� ��T�^o�������>e�OYW� *�'D�"-΋ $��(��D�R�5�S��j�.@	�����E��(ɸ�)��s�Z=��'�J����P��<Ȉ*@TT3���$O�G��`�D[�%�A1�*�(E#�����EXB�17�AX*��F-0;������@�G�|�`9>��-�C^+�V����^\?�7O/���c�xb.�ƍ��q���x�~į^Ǚ��p��r\��/oƑ�kp��f\�}7�:�˷�G��6�]�%k{�3R���"d� 0��Q���r�[�\b`i�PK�G��6��Ꮀ
s�%�"������U�3,�]`�!�*�։^�I�m��S|�H�tN�KF\3������"� ��iH��FZe2�
��Z��v��_��uè_3��m+���6�?�kO��҃�1�}5��߄m�`ϵS�w�^?��7���s8r��_;�������s8}�,N\<��g���ك8zz?�ڋ݇�a|��޴#��=܆��l�FW�c�N�.n� L��YL?�+�����Ğӛ����<��(���ǁ��8ra����.��ы������w�|�&�����Q��
T�/� J���U�!=BK
_��\����d�}>y����˹�m����g�V=Oq�����g����B3_�E���	� ����H�/��(l$�q��S�8��� �c����R4ڭh#Se��R�t3�st�T�tkf��<�!a�v���ꑸ�]�V�k�B�{�"��?�D��b�2�z����0<��������y���g�8u����.ChW6�8���1�@�|��s9�0m̀IO7v`�/���bףk���El�q
�/é��p�����k���}�yx�G`���<��t��0�譯�G�)O�mC:�5�p|X�%}��/�G�}�&֞؃�MH��8�O%�~��_��sb)b蜚��W�����{��W޾�����)J���D�tVe� P��`(�A��
	�@y5��q��M��\�y����S��bm��3�T���Ha�n�<oB�;�2�aIq-��K#�>R�Ґӓ�ґ"�,�Da��<]��s���q�>=���K���2��YB�˱��u��X~y-��r�K�1rt!�b��B��~B� O�b��C�\���]T@�:Ѓ��]h't5ss�m���ބ*�w�߷�}裂z��vB�y[���~3�� Z��P
���
�?���2��QN ���F�{q(�� �8x�[����� �j@�t_���<<r(��k@۸��N��	��~t@��=�"������%zO.���ŕ~i9�]߀�w��ȓ3X}y2��9����pM�V(�s������4$�e 5;�i�������}}���hx���������5������I �_`C�����B��Ԡ}h>�����._���ZX�{ &#/��-;p��E�=s���Ɠ�����`x�8j�b�9ݵ���AL]:"k�S��zApO�rGJ �#\��d )m�z^F�]ڄ��}�|� ~vV^߂=��c�{'�睃9��>/�M�(�Z������#4Ý�TԜ��~�S#��䁇���}����m?tt� V_��a၈���ZQ��	�K+���B�- |2@y"躟 �}>+�V�j�uj�8��U�X^�1��\?,$����R�З��?�P�S<���8gTS��2����({dB��p�Fă=m~�iH 5��	a���c��@����%x2@��g��Qa�"m�"�2D�i7{-�Z̆��&4fC� �LU"�*D� U�?��,����)�@���@���!t�k/�q�S�M[��L �#l�1Bi)#�s&��<�2<�'�~rS�B$4�%0IL���@�υ�8���ץXC&��i��vI�H�>)��@�p�Щ�T@)= �N�)d��,��`�DB(T%�ꉄ�d'!�1'�s��a�Y�}Ԧ��XG(�Y@��f	-�v�94��=�^s��Sz���=0�0{���ЖzZW�c��|x�/����[���M�vf%._�3G�؁a�8B@}i._ތ�&p�����Y���5\�u�Noƺ��ǂ�jԵ�
��#"��qNp���!�#���-���p�p�k�;������o�$x�9�N�d?���S�ʣ˥�δ�/�я�GF0<2C��
����#�8���j*FNs-K��^���N�@�W�jY/��u���@6�w���ct���^���kзu9l_��gwbÙXud֟؊��1A�zj'��څm�w`�ѭ8p��Z����c����vl#6�_�e�b���B���՝X�wVl����&t.����#�yv�Y��g7���m8��N�����Woµ;Gq���~���y/�~����o���<� �ִ4�e^P� �F@b�:I؜(�A*$� � ia�[Qx�!��f (�r:@%	�R�̩at28y�}=�bd�� �ٜ���)ο PYF2߇��*�M��N��|Hoʇ��<�!�y�S�@�>�bH�OT��gp�j:E�dx�G�����V�B�T�V)4�U恈��c׀��JX��Ý
�T��9;�������z|D� ����4�@>B���Tx��:�f���0��򢿙�}Q�?�k?9����~��q��+�ڰq��p[P��Xr�����x�����'��{/#s�0l�Ka2V�e��X׀�݃��܃p����"a�����w��������?���|���ˡ�A��|l�v�����-n�.����s]l3`ٔ��R�ߍ�o���q�������~��Va��x�w��o�£�>���0?����Xw�����k�`���p�L�z�7�R�S� ��h�V�C�:*�aP*�R�fS�0���'�<���O�⭃�r� Νߎ���\���H@����LXfxã8�Q��Ars
r{�Q�����C��|ck����sc�EX~�Psa)�j0�����9pt��b��(����ѷ�и�m�:�B��.�Zϱ�8Ѕ^�S׾�|:v��sO;�i?N��t��v*���l!l��k{7�`��m�:�4цƉV�:k���PI�wZ��@�T>�6�P!����Z�m���y|hf����2@+w5	��t,�Z���is[���|�kDk<\�F �������� @ �>�K!��וK��E!t.~y_[����1ry��;��ǰ��zT�j�OA(,����/B\\Q&���&�#=-�aa��5�e|F�����	�zƈ��Ǖ�ױ� �G����E@P"b␐��̼䗗�st�^���/�Œ��92������u�`t�z��؆E��X�k#���'tv�������ABS}>�\��0�������D�*�X�a��$4%�؄ڡk|v�z ���R��R���w�����0��n�Z�:���:��jD��*z?jf(�-����}����`>� ����C�i����,��>�]{��y@�(7��f�<h�k@s�#{1����!oE�0K�Z
Tp�(�VӋ��0�	��Y>�J�@O�7��ݴ�H�@s���X뀚;TDZ�4���PJV�5�	��ДI�r-h��1�	�1���6!��G4����O�g �	!�>�� �E��P_��ێb?��tՅ���V���#���V���T�r�Pe�Y��6׆r����)/D4:���kP��熑�|&�ə�h&��M�,ǘ�<�� j�@e9V�H>e�)6����D ��O��5��>�r�'�#C�A�x�[)@y�!9}!�'Gzr�[)?�>�� h(@�s�J<���G���x�(�:���EP�ӓG�e�1@���Ќ�g�9|RdR�����u���N�z�'�ק�^��)�� #� ��3d��0���\�<?)G� �@ UJ��2T� ��5�I�Q���A� ���5�џ�m��2H�jQ�Ј �F�@��ӵhGY@;���t1���\w4t�c|�;'j�}u9v�����&��Ӈq���wt���~�::��V���8sf5N�]�ǖb˞a�<�N�ǶC˰n;�W����N�U��+B^c2�k�Y�x8FZ�5���x}|�ɘ]"]�Dq�v�}�l��a��D�g�7�S�`���T_8���1���M��U���$ϧ1�s��:d�DV <�#�_�@?��.��_y"�r��]���6d"�%a-y��(B|o�{ʐ:T��&���~x":r�N�+�
��=�Ƞ�7V�́
Ķd#�&��YH�.BZg�jb�@����J4� .��Eh�ԉ�E�ȧ�%�Va��Ũ-CFk*:7�c��[0qi[i���^��w��:��K����,-��"��y\��
.P.~yg�j�B=���Pꉄ47��Qp��-�S��I�ZH�%g�n�(�rˑ�D�0F���LI{.:	�S#Ma,�0.'Q������~OH{Q��#�� �B��R<5
O�"�˷�mS#�#q3[
�|r-�4�MjAq��7@���kE��E����ɘ䁅x���y
PZ��=E��:#U�GPF���K�� epNoS��	��R�M�3Fm{4vT<+D��r֎J��Y=�nB�X�Up�d��Â+�ѽ}篟&u��)@�A.�#n�ʵ������#���������o�}g��D��ߐ������|���N�jC��f�,��7�.�ŭ�|�G���|�6�8��5]pYV�5��[\͞dh��BwA�u&A�%�T.K\X��o_�ۿ����=����h$��#��W[n�ś�<�xy���ٻ>�p�s�YG�([G���Q�}Q����?~�O��������)\y�n?yo~�.����Y���±��.��[_=�����#[`��y��0��nC���@�&J5�P�
�b�T2�0/��K��\u����Gp��Q�ta7�M#2+ �E��lJ�Ou$\J��P�K*Zex��,!ձ��DbK�{3�L�ZJ�=k�,��+���UXxbO�`���=>��#�:2D�c��0�	��`?Hۻvw�m�
�]	����}�9� =��s���oE;�����׃*��nk�A���݉Ν�h�܌����o7a�-[;д�]H�f*�B��5�PE������G��� t{Ĉ3 ��p7���ђ�<�n�VW�lS#���8E�>5��h%�6��@���O�E �N1@�ր֋B ��i)��V��I�axr�(��[��Q�m�׬�`7���� ���9J��� ���tz���������0ti)F.-�إ�Xu}�?>��Q���%�0�q����sS�VU���|E�!08 ~>^��򄟇;b#��_¨��b�c��o�ܩ��D !4<<�1�MJBVA
�Gmh�����8y�2�޼���k0�nZ��6:�����X:�����FB#���<[Kݔ���tU'��2�yT��r�}�/l#=`�ge�YB�'��1��G��C�p}V]݂կlŉ/.cߓSXs{+�>��&���W	���P������Oz�gH����D� ��A���#(ET��F�o�w�}R�>�t̺	�����ҳkE5����p��w���Y��YK�5V�����[VJ ��n��PQ�*��N6�%�r�jn�K ��n(	���!��,�9>���Fw�:�\њ��$�S��.���^c��c��"?��!��D6!4��l!4�M�7C��	�|��e�8J����O�x � N��e��B�D�A)��'�q.����\��kR���V��:p����0�S��<Ehj)Bc�2ԴԠ:O�:�:�g�( ���ZT(�P�%�RAW�g�a)�s���|6�Qo�G�Pya4ܩ�����Y��H�k<�C/L�b6[�VΒ#B���z2O�V)����V�^��~�<튌a��)�5��V��95�^��[�>�K_
���[��R�ߓCsj��`ß�j���z�$�#��h�|�B�!�S���h�?/�Ʉ�i�c`���$T��C�͟i��uZ$���) ��'�4%c	��,C��%G6�
)�PNs�j�(�R]1'��inФ�Y�й)���恹�.�Ns��t�/�*tL:���D<���P1�&}��i��<;6��=
umQhl�Fsk4��c�ٓ���T���{0��K�pe�V�bxy%�嶡\�v���-�N��(m�Cak<«� Q���`x��=��I�T'X���,�&��i�k�R�í�f�9����^�l0��<���M�֎�ǜ8[Q�MN���V�+˙�d�d̡s�Z���Ɏ�C�=;��(�y�tg�ɤ�3���]���9�rM
_����L=-�:^WN��*�jt[�d{��k��9�eYz�%B� oU��+('��J���c����Z�0.�aY��tmO�ku4l����ѺoK
<���є ��T�f#l� �#E�G�@Bd#| �#��+�oo:l��a��h�E@�;���Z��H<��%:$�vK�ZL���%ɐ\�"��őZ�};'��2
/��J賑% ��	�P��gF�������b�����Q�C0㥸�qj�}v2<Z����N14��iT���n3��O!KP�T��A刯��׀R�	��uQ��?;j۪��o�)��VCs[���aގ��j��Z��F��^,8�k����w�&��F�%��?k\���M���æcΉ����Z�u?/�#|`Qba�/
u���;������kWѴ�	�����˪ະ��w���ǻ��|xݛ�!��c�pZS�U�0_^
�Ue��TcZڮ��}�#�`�[�p�7�/��}���1?;��Xy� ^��	���<���+�Ғ��\��º?�}�����{�1|��~�!���]�x�>^y���u�>���ｃ�����,;�w�)���C�����|u9���9�ј��Yu�P(�|e �1�*H��R��v��N\��������p��i�|�&v.Gry�0bzPMB�޵Qp-�M��0e�7���F#�����H�P6�WU`)�r��Q���!\b���\�E'	6�������c�� 	��]��в����ʹ���$�����}7Arg:w��yK� �nnV��-�:��Ϥ��@ m x���u��	*�S�i_WCp���l�6�p9�(�<˴��E��twk;j(�[�PN�-#�NM)�`C�P_D����xi)F_^�����B��g5�n�0HP��.T���F�n�'�r�'�A�VAa�p�LO�Q��AX���l;t<Zo=D�?ҏ��B�	��<׀N���>������� �Oc��(��.��eX��VL�q k_݃�=֞�t��D �0I����Dx||�����Ą$'������npwt���#\��hn/'WD��#16I�	�)�CqM92���N�[؅�ucX�c-����iz�/B��lCe?�w����*Dr��6e ��~�S�[� �J���­(�����󆋯��� 3WAlH�QY݅Xzz��ه��&���Vlzk~z
�>?��w&�y|� �L���
�vK�5�r{����b=��z�wp�J;mo%��gas��7���!���I�z�M��$�Q*�����B��&گ	��9��\���&�>�`��*,8�zи���󁶢dY5r<�� y	�y+�Q��yk�P�N4K��jT��>i���5��MbMA0V�bM~�S����c(��Y\�n*趧��9��T�m�B\M�5�CMPl��P�Z"?�
���"��PS�|���yF�4ύt�C��"���糃�*@�3�����wЅ���l�ag>�j�7O	�胠6G	�Z�� �)�L�����$@y�P!�P�Ѿ��?#��td�g�� @y�O����T+���@e&��Ka�R.�vFlΔT� ��ҧ �H'ZC�~�%�9H
5��O�&�L��	<J�Tg���B#����yY^Х��LO�%��M%<%�B;�s2�Yn"l�fSf��Q�4�w�Ch�M���=XF�2\6��p�0�K�ܣM�C���V��p�1�}�ab �CX�{bm[zܶ�,z/�B��� ]���עm�0;�XX��9�>Ύ2�J�)�)J�0ȇ·�L�U��c!J���4Y9�o�~��?]��M!�ʙ��T;(��C1��P�m\{��zo$�D�β�L]��$,�� ��Hq�D�$R�}�%o��s�l�3݆��v�ˮ�Ȱ�$݇v}fW�er��R��B7��9C*�^t,�%O2�%}�&��lI���+g8
�W�?e$J�)݆>7t[�t�L��j��s$IKyz\�y.�Ȳ���c-��K[t�B~(rCq�����OQD#���N� Д����ZR��p{�1r&��Qm��&\�����N^�}�So'ο��9C�G~���E�T��>��m�enR;Q��3C��+o.{.?��;ka��[k�vx��`����ͯ���5������_�����
�g�x��`E��p�g��oR�\��WZ�����<Ģ�����K����*a?X��+���_�����/=���5��τug6�Wa��2X8�'a1� Õe�_S��[܈]��D| O@���;�>���E��u0&��զa��q����o?����{���1���0+��htb`ߜJ؀_=�����ￅЋ�o��G�p��X�s=��#a��eg���o�z�����x@�
"�ה����D@�, ����h���K�͇j�%��6���p��Q��� �W(;��A|q��L�e	�l�T����
��Ap(� P������/*@�6��D7�V=���]4�N,Ģc�:�s*@x ��0����[Zд���&�ܲ�pIm��N����"�v�r:>9�F
C�b����������J�@�v:!��n?@�"��;�wf^Y����ur�'�r߾}h:L�8�M %�8�3�z���w�CeU^��5B�5$�v4N/�(�wѥ���<Lp羳��x���F��.���v!��E=��ӌ�%<�˯N`���������@�������"T�7 5/fVp'pfgf"=%�NN�05���-,M�|2����quCLx8�"�����|�U!��9�(��`A򺪐�D�iY�K�%%����Hm)@|c:�(����J�_i��B��;�EV �c=`�ce=H(H@b��	������	zp�n�ƚW�b���p��s��`/_[-4��׹|k�� J��z5��5�:���[G��:$_f�
 ��zs:>95�S^2@9�F>� ���@�
��zj��/�	��=�]ߎ�u�&��.&�.��B�,F�2�>��|cJ�).-+7��w�F4�L_,��Ʋ,_!�ҽ0F���p�2�П��4wtB;�]О������p���ϧ �� j�@����!���w�E��>"<��OZFF�w
D��&��(��K���W�y��#u��)c��� Qu-EQ�ЧMl��S��T��dx�� �b��z�B�����Wu���zuћ����ޫ@���{	ћ@� ���w�6���8q&�$N��L&ɤ������fK8�$�s��k����^�JZ�_�G�}"�� �- 	DiJ+�;e[���HO��Xy�t��Q�@(cA`�j���BM���b�n$l7N���=`ܶN��:��q�:��c@�<xm�
7�|�H��U����_�A3�y<\֌��)����*�~�'�=���<?����Tw�L�^S=�9���g5`�`]�<�[��Xw�Ѝ�������<�/z��s/~�D����p���\�8N����ѓ�ǅ�Kns�g&�|�vĥ��O��7�����|_�����3�=n"M��g#!�,7��9�f�L�L iN��s�b+�?����	��PF��׭�'�:b2l"��X�v8�#�u��q0�cd{
�'p{�¦�2t2,B&�G�<�;��{`=��&��k盬�c��b,%�x��ȶU�$�9DO�m�4��L�M,7�	3a�4����Y*v�=����)}>�3��6k��Æ1˙��+U�+U�\�>�
��Y��{p�Mq�r�P��/uh��8%�����@�ߧĎ�S %���%�*l
���?K��H���W*�ͮ�~3�
*�� S_��
$*���M��jC� B�4N]�� �s2B1�2�g�QԺ%�v��+7��_�;��'���$���H�կ�'ct���Y�?��O�ϟ%|N�����/�ݽ��ù�t"��S1�0xn8^(C��V�����O>���}�>~�]W1>;@Aq��;����\��\�;��br�V�Ԅ{����Ⱦ��ϐv�Â�br�y������Ͽ����C��¨��蛽	���AP��SVc}y&j޸�����<���_����Ƌ��G?��?Y��1l�BX?Eux���[?����6�cC��~�X�m��sa�}�C��:h&l���i�d����%�8x�g_���W�q��sx���xDL�6�2"�c��x���9��8}7����S1�����wmV�,!@��5	@�Qv&yģ�3�h�~�R�,=_���'��l�A�4AR�̥$�����'�m�R �<���Oh�K��R��+�����G��N`���("C����9���]�Bx��V�=���R�=@��xR��E(#���~�"��M����Px���$|o�G��2OA��S���є�,5Rqƹ�Ь�\��6W+:'��]�y���ڀ��P�V�t�"�PZ_�����aI��E\<�kHV-]�y3�`��٘=s:֯^��m[�~�
,�=�̂��&�d$#57�	X��c7�X��+b6aY�z,�\��k�8z=��oƒ8�v�G��ܰ��S����31n��QK��w�Q��k}==���p6�[q��Wp��8��Խ}uﵢ��f�_��7Ag��r�9����{��T��q���Z?����ݐ����(�Ǟ��OIL}�Z
>c	UYO$b�h|cb��=&@�Qz�r[v4W�z0[v¿�xW C!*�����nG(���<���X"*cU�(B�1@7N%B��e�I(�z	�w1�&����ܵ㑽f�V�EҒ��=� %B��"4`�Pt(����s����j�@�?�&���D��\<�%H�
��' ���B�Q5�[�S3�i�{a
3iDo��Qװ�=ѿ�3��mы_Go"T(r$D�P�n�*��vy�tͧ���JT�������f�2Ȑx�K}[��{#6��q]5�U�C�<�=s�̌�ɜȲ �d����అ��:	Λ��q�X��<�;f�/��O �?��x̺�pZ=��N�w�4��w'����2^[�N���0�����i��>�M�w�D�����z���}��<���<�gc@�,���3�����X����qZ7J5=�_;��|x=�m��>.|Λ��v��9�Hc�fU�p�}�6T��3R}k�
�}S���P��	NbӒ�4#4Ͷp�?���������l8fD�Y���$��'�L"��&h범m�[DM�e�XDN6� �ܞ
��鰍����mFd:&��։Zަ��D�z��2f*,�	�P�aC\��M�y��I��,i�Sf�,�I����0Ϙ���\������]�b�� ��=i�{���S�\��O,.�e�
�s�KV�v�ZX����.�S��Stm7yO�͍�f��nz��4��7 ԡ�3�^�J�)R�+J �ic4Ƕ��`C:>���Qp�q
�r{�����L�4�;�΀Qǚ�����vk�g�oS��ň�H,�Mֵ#�uz�����n�׿�7J�5�i���=:>%R��V��ǴO��g�G��=��G�/��O��7_AV�>�=��e�٘R���ǣ0�p&�E��z\�Ỹ��[��Ͽ�W�o���ϰ�h��l@���p/�Wi ������Z�-��Qt�	mo�í��;?���GHn/�Р%����_~�@�g``�6����r$�wm��� l��C��Z�{�E���-����ռ�������!��7̓��i�:s���<���x�7����]��9#�`9��_g���|�[<f��3�5�Â�"7u�^�K��.^��.�q�	�{���G�P�t���������p]6�2�؂~pX<}6�ø�y��sbaY�*l����]�8ry
Nf"�M#%��}*y�s�ג�\.s�N�i�4�m"~x���T e��8^h�R��4d(|��i M�zRC�B3!s��} �E0���6�)IDp|c"�
�h���8�d�����]-A��<55��7����7�L��gpml�JT� #PU�S��KZ�1@�/�B�%C܎B��ә� Mo�Er�/8��O�f��T��d򹤝�inr��^D��ǁ�2-�)4�yGo�ī?x/��U�������~�G����h?Պs�[Qu�j+O���a��Y���v����9�Lc��84t+����X��\FȆ.ǜ�e�%	_���T;'o��I[�b�9v��Y6��D��0�$:����\Gy`u�?�]8�˟���}m]E=1]�F3��:�*�sϽcH��"M�����1���F�z�XCsg郛�V��Қ��3y*�Լ����%�O���4����Ќ�V@N&�����3���w�Ń�9]�	��و<���=�T���>%�GBUS[���`n�>�VeRУ�q�6n���[f�l�T�����k�D�d��L@S�z<�V�CΊ1H^�"f��"t��AD�`��sc��� : ˧��Rt�x/��E25�ԾX�}˦�D�T?�uA*�q��@g3sF�#�0}xOL�p}�0W��c��Q��N��'����Nőq�q��/*Mn��� �&�����.��>���� U�M�XIU�����c гFo�i���a[5�����k��������'K��j�(�n����i	O��S�3`*z�����x�I<�m�/�ԃ�t {�x{=w���?	�;���
�:�`��aQ�0,r�7LT�x�n�	��S�a|6N��ҟ�{�d�n�
?��������	��mӈ\އ u�1����ǎĨ<?�3��h�r�#/46����1p`lV=[��J�Y��v��ξ��� 8�6rߦQ�:#UO����	����M\���u�0':�w��9�i4�� "T2N��<b���.�䶅T<�mItJd�U$ʥ��<��	��p�7E������$j&�L"Tn3����Ħ�i;M-�⦫u�T2�bxl�4�%�ɂP4� �T�u�,� ���`�B��.�y���\��S�Y������l��,�e�
O�}��C�)[��D����&�2��aOmd�m�T�1�k���e��U��P��#���J�	@�J�hMs�u�8��)�4���;���2АI���\�aPc,FUF`mK6�o���P�r�_��_��'%�m�!M��B������4���50�O|R\�Η����C�ߟ���S1�z�y�>�y�*c��cSs)�~	W��^��gx��p��wp�����<�����;�q+a�}f�I��_}�&V���/y�x������q�w,���U(�Ѥ0��O��;�y9-嘔�!��)��=��f�	D���
kJp���1���|�׿�!�������E��:ټ ���#��~�)�}�n�� ���!� ߗ��;���wa��|DU���fԾ؁��^ǋ�?�˟���>{�+ߺ��/�ŕ{gq��yԝ)Ǫ�U�l�;=�+ŲA���o�^�ſ	���b*�6͋_�婫�s;3��;q��>dT%!U��9I\֧#�&���L����d��R�ҙ4�S*K���7��*h\U"�P�'�pe0!=�4�.�k Jh)�>���# t,V4���8�O�f?@cUS��3�ȹ�B$�L&8��ͩ� M� ��&.��z�A��O��g��y�WJPtu7r/�Y�;)M>�a�S�)��t�Z	��)H�J�y�B2:���jꖜ��(�j���8|�G�T�حj�8������~�?�w�ß��������7����������O��O�}|������?��p��u�*)A`XVnڈ���`���8�-Ĝm\߾ 3`f�"L^����b��L�@=�v*�_=C����p�ke+X�Z����?����{�������o_G��p�^5��x\�Zpu/��Fz{���j'�;�Dd4�f�PG���#��{�~��H��i hR!H�J�3�>UE֟Pg�I���B/S@w���%H��'[��������E�@��� t$LU<�*c��K"&�p}@��}5�����X�[f��P�f2JWMD���عbvr�k��\5�+ǡ����c��tRG���X8!�`ǜA�Fpn��k��aʹ�X%МL\N�Q�=���d��~X1}�j�+}@e�P�'�R�4��S5�|2�O�笑n*���2��IH��S��Dd��>�Gy`�x�sBo?�x����
v/;"�6�N��%>U�f��Ө6�M�K�2���V�Vb�m�� jCx� 0��n�d�O[�S"S�@��e�)�E�^���GF���o�����o3bԌ��o5��D��k ���+��*��&c=�VF�Z��%�)Q ẻPs5�6��"2������2R�DF�U��2Vk���ߎ�Z� TMb�"U6��i̻���ǒ�=�M#5\Dz�PFO�X�� �,7����`�e��	�m`�i,��M�[�L�b�L��iG`
�ܶMA/�'!h�n$d ��B� ��2�D��л~���ބ��)����qp�2^ۧ��
�M��6}�M��iD�Tx2n<��T?y~Wƅ�O�����:o�
�-����p�c���'�i�ǰ�s�&>m�������_�� ���ָ����"�z�%���K��!�A�U,i>+�%2	L=PA�E��̙�5R5��ӑi��Q��u�X1��i�|
D��y�U�4Ϙ��y0�bd`!	!*5#B�Ì1/\���� D-��s{�Wºd-l�l�=�hå%AjΘ���Y�BS��|z,�4*��)�1>��5Q�4�
,�d���N@�mki���Rǧ4����.[��������X;��D��g�?��a��GΣ (�4��z����҉I	�WDM�S���8�<���I\�Mi�&�A�a\"���j�i��g�t�tj،��:	�YW�gCz7����l���I#�r�oC,V�c|]6���n*�5���
Wo���~������~O0ʐD2����򯄩 Oں*�1�j1�����?���g�����������gO!�p֝��ĊD��F�z����R����7�<�W�p�;���Oq��7��w�Ǐ�k|�ǟ������Q��k'P�k�g!�|���_��_��~�w����{��^C`}	&�m����Hk=�W~�9>���җ��l%�$o�����/�w�6b��wm�w�
L�ڎ�wn���w�7��W?�^��[(�P����b
�N���>ƽw_��G���O�������}���'��~������?���>V��\���\p/~�>:޼�ӷO���f�}pmWNbC�F�_2��[�s��yzl�߸�#�ſ%C�fbB�|̎Y���k��x;"G���{:x1L���i�^/����,�S	�0�:UE�S	HA����f����~�zU�>MN�T��@���쬊6J���D\���(/��d] �7ɍ"D�N���t,atxu��~<"��q�	n\�[K�B�4��w)D�s1J0Ϲ�<Z@$�H�L�4��.d_.~b��SD����󹞦��F�����z�iP=�7�����P������V�)�x)W�J%@����TCU�������v�M�眅��� F�j�u��WK��](�} G�^%�nU��rn�u���?��_�󷌌����?~w������ǿ���DU-f�[��O���1j�H�Y<��L�d�g҆i�v2����F�g�`x��	~0`3_K��Y����[<
����S�K_���_���~����eԾ׊C�Vc��C(�y E7�!��ξ���w.��r@��, ���'��]Ve -&�4��$5�;לmX��=���.�Ԫ�R���}ʶ1DF��f~�Zyi�}*��5��"F�	n���w��<��d�+���@��DUݼs6��ʖ� "T����A��k��#�*�����q<h	o��}�f�t�������粱ع\2��b�`��.����#�R¢�C�F.�P~`AD�����D|n������)~X1��$<�N��q�/VN�UD����r���ԫ��)1n����� j@�lbs�!@{a��G�Ą���+&p}<�8C��~\��c���prg<�*Mr��NgB�������V
��
�R��g�i�^<V�%D'c!K�|�� ��RL#M;����+�� G0$ؔ��B�T��R���]B`��\s�hXm!@���v�x�o�@�N�s�T��̀K0q�c*zH%t���nĥTF��Gܙt�:n�g�u�[��ӞD�ʖ�p%@�	@��骊��q
\xn{�Յ����9�8�!���s��O��f�����<&�83N*���pdQ{B�ޟ�d�N��V"�(�!Hm6O����k�u����u���
�Ƞ@V۴H�N=���ܟ�&yAkn�'�կ�\O��|Vk��SE���y��o�)]"�n-������용0cd�B*�ħE����� P3��f��V����l�3g�s���%��d)�
���g�rXI��b��ZŪt-���+|ZqiQ��R	5���M]�w#���^�$@;">���Sz���DA���}RUUP�����&@U�Q��HsZ.ut��_������m�oy<�6CES���d���@�1��ap�Q�����(�0 �g}��nJx������Fb`m�6'a��b�x'nբ�B%��<��_�����������O�Acj �ӟe�\^9
 ŀ��	P�ʨ��>�����~���@��vD�eb�L,��Ĩ�D���A_�?߇���N�8�(}x/�۷��ǟ�������~���9��ŗx����������~�s��?��_�����G��wx���j,ˋƬ�1��cR� �Z^��������m�Wbd�z�ڂ��;�wO |v�ót+�x�蛿	#�!�� ��_@���x�����O����1r�N��Z��_9;/�������'x��w���?���C|����
�������?�G��|��/���)����_��{�����>���[�p��kx�ݻ�p����O.����c�&N�#��9��JgX�\��X�Y1˰"c��#�h,�N��L!�/� 4�ɲl
B%)5DS	A��3��O�(�Io�R|�8�ui��u 5N
�)P���|��*�|\-�/Q�6@	I����Ȯ ��E��A�d "�~��D�t�	 ��OFHM9�O��T ;\D��"���jJBA#�?S;�E�J�3��kHT�P� 4�(}@e)�4I�xS��$ӵ�& ������1�R]KU M%~���'<������$�r�Mֹ�����l��|�^�G�콻��ۇq��>[��w����o��#������ٔ�U"-,�fi?��߷?� w������^4Bo.{�ו�pz����{�|�=���f�zL���q:�ǭ��pĝ�B��F\��m���C\��=�~�:?;��wP��>��D�n��؍���!��i�uR{6�
M�&�%[�B�!4^��4TA�$��mҬ�x%B8����5�I�wY�OI�9S5��$�R�x
F�z�[��	��O��W�LB<��7Q���BQ�^�ݧ �xB *%����! �
[��Kqp�\�Y?{�LF�ʉ(Y6�KǨB�W�C.培`�J�$/�ą�!n�0D��&x�@���3bˌ�h?���+e�t�D?�\9��L�5P��EpJ��H��P���:B;#2��S3�"��D�P��2�9�0�#�s�������	n6pq�EO8z9u�*ӳt���� �����P���?��l��f�`XK�����)� T�G��P���Y#�x�@8�*�sJ?E�Oƌ�4�(#�>���jI��(�6���6�@���qp��`b����Q��E�4�\:���gG@�r�w�����*8���@oi6K���D��E�E\:�~��S��񱜸^���D���1{q�k�48�R�u����$��C���1�����!nU�O��!��:�����1N�"�q,ƪXH�ZF�uJ�Z��i�8���L��S"����%�(��g	��%:8�b��M�&@�z�t���蓼��:<Ւ1h#��#:�N�g�2-��a!�$>m�W2�`]�NŊ�ܭł1c��{���O�&���B����'�)�|
>%ּM�)sn
8�mo�V��J��*@Q8�T�&H��o�i }�h 5n~�Gp)�k��5��� U�o���@|6Ƣ��4��	@�z1���1�����
���*T�X��K'p��)\}��޿�/������x����#~˥TE�|��L���2ߊ��c������7���[�T��%�X\��ח�������~�q����/3�r�Fbؾpl�Eܞ�/���wq��7q��7��_>ė��)~����'�~����|ݿd>�����Ps�o�b�l�Y�狂�|�5�gֽSx������'(�ބa1k�/c#����� x���}�Vx�mS�W�#r�c��${�<>�ݿ�+^�?��� ��q�n�����Y���?����O��?�K��+��ǅw^��{p�͗p��m\y�&.߻��/]ŋo���s�Ue��q.慯@��f<�����5�~tA�a�Y<�7��{�~�L�߹���3~�s0<r!&D-����X��	�Cy��T�.��K�HBBE2ᙅ��lb���LQے�Zb� T���R���`D2�DP*���P�]��;�6h�OOþdF�)���lJd4\mj^�K3\�Shp� T�TE��`S�S�/�SMr���;���C�`F��Hj��P� �s����U4�?��ͩ�_���F�y@y�2���u���>S|Jd��gR�V���(��8�ϡ=_U:�z"kx��8Q�-��J��Ar;�����Q�ĞN�\�$�i��y%��PtkJn�F��2T�V��������R-�~�U������=��?ş����]�_�)��'���[�^BpJf�[���G`��a�7k0����\��e&Ǯ����C�d�,ŉ���ԇ�p��;h��&Z>��K?|��z-_^E�-8�V=J_>Jx�!��.�^�"�r��"�˴�yH����Nl��T����D0j���d�#�M��	����[������,���Nj�O�g�t�gt]2�j�<�HE��4��|�O�oL@,���H��E"�ۅ�{P|� 2�w*�FMSMp����>�@��W���]���pp�\�0��LQUP�gђP�e�����yd���!m�0���L�����7�L���2g���n%2�N�Փ�aդ�*�'�S۲T�&���iZ�s@�q����j�;f<�AtJ��Lg�T�G�a":����\UK���������᧏��aO�:���^=�n�)����a�T>���*��T��Ml�O�S �*�� T�C�>%�a|�]��ݢr3��F^�
Q�c%ڈ��c&@%4Mc�X���l�}<lwL$�&�z�$8��@��Y��t�o*vo۹� u����TF�m��%�b�#b.�:nOB�;|��G�l�]�>�K�4��
{�!b6#��1|6z���q���U��Q��1=��)���2$?#s��3v<�Ğ���9F���3��a<AŚ�Ԛ����?����>���p&�9���c��� e�����c�̯�7h� �$P��'���C��i��t�S��u����ȶ��,x.��N�
s5��*��v;�����,]Ɯ1ۭŜ��
�ޜ�|��.��'����(#ۖ�	Oc|�v̧����j'�e���vV?%(�� �'�$v�>�'��F��c̿��T�4O�S�܇��B�'_����zs\���Tovk�@]O�gO�'�U�k����}���w����T<F4�bF/�/c��r�ݯƅG�q�~|p���|���◿�1~��_����Gm�?����T���|�����wp�L%�w'cEY,�W�b��4<ה�����A5Lm<��LF���u�#�q0
��y��q_��	�O~�c|��?�G_}�}������c����?Ç��1j\A��,(�Ǥ=�T��Eb��P,ڎ��ո�_�����o��8��cr�?ߟ�����ط��n�[�w;<wn�[�*�؊Ď
\��{��Oq�;� �e��,�_�2liډ��\A�7Q}��;��}�0��E��j�U ��
NFN��V�"�<�G�}<��6�y��m���[�g���q]����Q�z\��K����tU�;�9ã�9�gŭ�Ҵ����v ��O@2A�B�%V�jЬ!H�x�]%�l}������V�wʜ�Y�JS\5��>ӛ�U0��T֥_ha�`��$���h�@]���Y���8��S��T��
8�;�� �H��hw ����
*��myȾ�9�wBF�M��Z�&���ij "�T9�R�T!<U�NhvP�U�*v���%����7�m�S�?�	nT�Tq�U�RMm#��s��,5"o�ۢ%� Mh��R�������e~^W�s��׊Qzs7��;����Ps�nř{����	�^;��ow�!������ѿ��w��n��"*�4`_[9ʯsy�Eg���~��?�C7kQ��,.|~��.���-����������Wp��ۨ���?�\F�G�8�z-J�<v�=������&C,�]!<��S�y�,���#�c��޵����:<���[���Afk!�� �9I��&��L��,�-�qR��ܤ0�7���KBx�|��i �}A%ZP�G*�	ѓ�Dm��~��2Qxn/��� ���#�������~��E�CM�T������8F��2�6LǞU��s�X���G!��Y4RU?S�E��AH�2��L�;�L<�}�s�!r�sgBfA����<}06N�u��c�$�������gQ���`�ľXA�J�P�B$S�H�Ks\bi�H/��L}��@{2���|OL�����=�Q/�0������ps�����'�p�����T�� U�$6�~��*�4����h�k�ʀϿ�OB�ihZn&(�DgW��>���?1)MD;�)�|2���}��r�8��j�$�M�s�l8��$�$RY$4�"J�:OC/bQ�2�H���D���;r>z�\��,�o�"�F-�����[��1��_���X]���D�,�D/�+�Lp�E.@�ȅp	�琹��|��9�x��yp��q��ׁv�sq"N��|�.ܯe�ږ��zæ�!���kU5L�&Ӗ<�l��=֌�-|���җS��)�Y������K�Ђ1�Ѣ�dF�~�u~m�!���&Q�p�u��~J\�[�O�e��W�|Z���a�6�saAxZ�&��`�� ��<����Z�N������Hs[��5p(^�bY�^��r���� �|����-
��T�)�!��<�V�)�Tslri�O�%����ܦ�Ķ�D	�:@U=�)>%���[y*@�(��$<�hUL�� T�iU����L��S�6M�=>%�P�F�n'�l">��>�<}	P���4���j"1�&
���Pr}7N>���G�x�[���7�ʷn��;7��{/᭏��o�����_����TE�y 5��w��>��S�ߏ�Y�XU�e����!|������=x����?Q�۔��8��Ģ��p��E'2�{�?���ׯ��k�p��ub�*^���_Ɖ7����W�}����[��`��G�y|��OY �]�� �jr��"�a7��bhY�˶���6���j���F��ڷ�{�^�~9[0��c��L�,K�����3��6�;c-����s)�1&~=�E�ƈ���υ/ǀ����?�Jf�w�t�o�ߧ5/�y@m��2�����3Pq��}�>��]�~�"v��w�h�����������w��C�4xG��0���@ώ_��I��&{J�y8��\����ޕi*RMpr��3��Pd��R��!��*�����)m�\�(c�O�P�H��#,�i� S����6���D����HT�O�6��x,ƀPS�W<�Mx���� DێE���2Qj{��VI�ۤ6A�������@��W�P5�*	:e�PQm�O�<e "}J���* �G��&���^|
JVi�Gx�J����a4�O\��`IĨ@4�|.���U.�!�R2.K��"^.ƾ�{Py���C����؃�/���*p�n%N�T�ƻ5��S���g���\��.��!ھ}-De�'�p��lx�2�����K�~��P���_>�#����7��ć�Q��e�>�C�+���Q��9���QD��]�A��dvd��~S��u��L�9"���9���6�yO�JM���6��L>E���И�" Mn���l$�*(����]=��u�Y��CDu��֫��)�)������>�9I���F��� }@�Qܱm{�p*�Dcsq 6�� ��^K���4�=�T�=�mm���Dhٺ)� D˴
h���\8iDf�A
�)s� y�`��Q��9C��p_Ԍ��1 A��YC@�n�6 �&��.���m��a��!h��冦�K��`��'�A}�`�/��¬��a��ў�9J����V��Jt
�5yDo5���{q�S�����P�s�Pw���!�\����^�p�9C�t�j�w{��0��p��ޯWgl�m-��
0	I�>��/o�R�Mc#��K,"�6�o�O���� /!2e�[�Se�(V�{v�SF�tZ�K��z8C|��=�2�%�?K�S*���V�~���8�(�Љ�Ps�N&8�\Z>�r�X
:<�N�L?X�":s�眾0�+!<�1D��|kP���Y�4�x
:�V�+%�`��kd�H����CxHEڨ5�5��wSk.���BѸߡi^�G��#���+J���x��X�v�mc����*`<�	P�`��I�J5�N��D�3��CA���6�ɺ�@4z|�W�3~	\�P�Z
D}㖢O�2��.A��q�/~����̍蓴���CA�4�%@�x��D����[��1�����=c�%�H��9Eχ�9F�vƖ����9JBpF�E���\΁��m�|�3T�"��)��/b;��O�c>�����ڼ��O��b��mMXZ�D�O��~���"F��S�
o{���&Q��ǜ�&�_�ę��$	<�<�g�<�s>�%Y�aA|Z�.�e�bX,��iNxJ̊%�`NxZ�Z+�f�Zؕ�c����n-
�e�j!����}�a����҂K�9aj&Mp����(�r�ږc��IBT�W4���iyDB|r)��2�.�X��)�<Z#*	8��Lc�uQsk��\�r>�oZeh
:<�j?(�!hC�)0vQ���o{J��yn�)8Mj/ �R��+�W���I}]�t��H0)�mٯ��)�	*�ky�Iz�	8�o�#�)�W?�4%�����4�ex��* �,��FM�h�G��#8�j-.�ٌko���7Zq�sx��������*��:�7�y��}����7ԀC}���b��?&7��RÔ���ǿ�p9�6���9�(�_����Ru�~���ꝫ�9��w'`^YfW�bA3�)}y��w*	}y��W5�M@_Ƨ!ލ	�"@�p}Pm�;����1�HfI�h�,���H����{"1�4waBI0&������?����x&.��@o�w�fxl����R��yA8`w �
���y�����O�����W8�ع����5a���)v!z���g�Fxn�K�J�$.���E�;��"������D�s(��ςK0�N���n& �'�!p��d�(�:����w���_����/c[N$<�� ��p�ÿo3`�Z�L������c��`&� y-V�l��]A��$"/���UDUA�eJ��3��$EAT�N�њ&K�M8H,�4�"�I;)��m^��_��[/�4�L�>i����Z��EFѕ�I*ђ�$�4��d���u&��� C�٭�~�"�&���_-�#e��(�����F�`5����,�\c�S�,�y$ۏF �&��!@���&���0�,a�F���!���8'�|D�{X�~?��=?I|r�@��Dft#���|�Ȝ���6��������*���S�}��MLWO���<eP"=�܎��x��h�Kٖu���'�k���Jd��g2�#G�4�|�������,\,��k%���o��ћ����u/Eë�Q��q�|T����q��� Z@����E���":�����"n�����C\���8��4}@x>j"<P�V�k�!b��ku�s�%������^�����|��Bd�� ��Lm���,��\�t�g�:�x�:���T?�Z�<�m&^F��Ⱥ��
<�������&��"��L6I�)�ܧ�y|�6	�����LTM?�����~>���$D���=oJF
�%񳏫�Ebm��/;;ʰ��>d�#�*q�����E�P�ͻ�u ���0;�;*��� %8�QUq�����x�^]� ZF�@�؎8�?GMϲ�L�V����㐯7Ý7��g�)Dg1ڙ��2q�@$����#���q�� �����?�/�N�m�bی��2}6L�5���1�X6�K	�%��q��?��_��>�;�/f���7�p�3�f��G����4�S*�
��פ�MpN&>'��1��m(A7����q@owk�7��ˑq�3���B���^Tpٛq'(�	�ް"@�J��ӡ�;����� �$
���vld��W6�.R���C�`�X�S�����w���0Pk�S�����2jz����+ް!>��N�)D���)���B|Z�$8%�� 5����|n��� jiP5����xJ�Ns�l��C`a�n�j���a�i���Sǧ��S*�F�������|Z:��[��thZo�����n�)�2�c�t���)rq6�Qsyq�.D��O�:q��$�d�`:��dw�Bd��jbr�������E�x�,�o�rf����&��N^��E�5��D�{�2��/" ������8>.{���;FυU/H�I�R"�vѳ�;�1�պM�L�
<��P�t����&�)Ĩ-Qg�sGMՠ)�$ e�q��O��g*̈�'b�H>s����Q�u��0#<�O���Z��Xd���E��12�������Vħe�2�8Mb�k5,�%kU�O�Z�S�q��ea�G�	�{5�Zج��s���ۨe���9H���D��aއ��+���8��K�x�J�5B!L����Y=Tp{���"ǚF�>Ye|Z�����ww���Ӟ�<��qO<u��8�un�'�%�1r����~��C5��8�(���d�X#��ܟ�m2��6�퓑�] �}
����iT�.�ߩD5�4K��g[2<Φ��\��5�Xߐ���|�} M�U�����)���sx���x������G��/��_����60�_�L6��d4�R�3bX������_�_������������?ɠ%<^�����_~����*:j�;k
"0�_���1�!�y�݇�}xaޗ�}y��ېDt&���۳!^�7/����З�[F�T�~��я��C,�oE�R�d�2�vmF��L�V����c��{4���}4��;/�z�۾mp%*]voAO.=�����8�ۉ�mp�1��nUq�C�r�;z�.��T�nśЋ���m�&��p)\���yka���Y�ᜱ=R��9i1��.~>���>����;:}fa��x���λ�q��E��J����蹙���1t>��M��)������B�L�_�i�*��h����uY�)OV M�p)Lb/��uҔ��\O P��y!o��	/�C�&�">��	��aqŤ��B
/�e`��:����Xy���"8�x�_Op�uIFpJ"����^�"��&��g��un'�����e`y4�
,#�r��y�&H2x,A�t��pD��ȹ��P+B��|$A�g�ݚJt&)ȥqQ���g,ᙀH�K��s��(�4��ei�)�8&4+�&nG�|�L�����4�U�O~�Uœ��m�O���4FCzZ��qP��ĵ��|��'4�����%BS�i�\ʹLd_)D��b]�E!S|)%WQvc'J����w����8��0��v���W�q�a%*^�Ʊ'p��Q���4|�$�?>�ӟ�����8����ً«;�}!����K�j�C�˾L����Z�Ҽ���}l�mg���樥l�z�@�-W%�lR�L��I���:���������x�2(�i-�g'�q���bO������}[ş�����}Je$�S�Ȯ/Dre&B�s��h;�mƦ�m���E[��h��*x����0�	�K���5����@E�2U=�G�������l��0M�*-\>VUA��P5�TC�P��M����9g��F���5;x��i�(#�~�����)��|���R�h1!���7��Fy`��~X9g���y����Uf3��
J��(��tҐ^�Ȍ����{a8ׇs}�����s���TA�Z�P'����������PkiZ�
[�rJ�ӀO�i���n����
�T�������Ԧ�	�ͣT4hv,5Tj�4������*�c� �ߊ4�57�Oc�:�N�c���$� �(�ΞD`��F�W�6{�=�<N�h��^D���=Cg�=��$.=P�����]D�JS��*�j�m�]0�3r���<����%KWh!jا#Ԗx����	M�p��On�}�-q���0�caʥs�,��9�6V�s�:B�@��1�!�R�|��*'��%O#|Z�́9c��7U�|PS|Z-�u�oP�O�z��N�}[`Kx��
ۃ��(ZMK�R�)�j�i����W��zE�$2ϥi�z)�r�&��+Y�����Yڥ���'`�5��k���0:��C�z~�D��idw��4��lK�SL����!�s��ǩV�]�2`��~y���UZD	M'�S�f����P��
�^�����+MS�PY�nM�w{*��R1�dF�Bz¡,/G/|r����K�q�ch�74ᵷ/�_}B"�4�:��jj�ȚPQ�*��2t�D���mO�0����'U�����������݋Ȭ*��ݱX�7
��cZm�5faĩL��v_^���u�F�}}y���x7$����DـP_"t /���?/��������,��e��/ӟx�,����߉0x�A���U�#!�f|��<N�uD@�;o�:D�t"T��@��� o����׾ ������Z�=���s�ږ�s�:�g��s��.����B�&/��$e��i�m�aQ��|������go��+אt�>+'�y����H�^���S�C��$@��b�4��؈�y[�qg �����TT�	��v�4�%H%�\O�m��������/�3�>C�S�)M��4BQ*0��d�ĸ��N�F?@Cx[Xu"���Զ��1��D�|r�T8*	� T�M�i#K��B�����D�T��ݓ�Y�Rƕ"�\�G����?{��2�`�$N��k�k�6
���AA ��ҿ3^�z�;.K}]p*UQ�� ��IF�����R	��RA��<��C8��5�ƶ���n3!u��G�J��x>�R�X��Y��q>i��U�;ґy!����wOڹ4d_�F�U�?|O�d�݋�#�3	�tW�Ko�b�K����^5�Q�]ȿZ�iܑ�T3�B./O�Ô ��i��SGh����c��NCd;Y�C&Y��J���9�	nK���<e0!՟�1qDe"� }=�]���$"�:�5���;* �g��#�S�תʟ%~�c]���x$�{��Z�⳻Qtz���D���Ŧ�X[�K��e�l���#;P�-@�N����E����f1�P�5+U3܊��8�UAB���ލ�Q�n2v���bi��b���
D�QqSfF� tZ?�OediH���3�#�	eBf`"h�@L���*�n��� ��U�5�2��0D�TAL�3�b3R_���'�#:g�f��t":~pOL�F��R ;�7^`F����Ĉa��:���N�pp������`�Ӄ �~��I-�����oS!�0���F�����}ak���V�Z)����e4����4�^��Q��rL':��~Lw���X1��I����ai4	�!S`J��&d:�������(ʶ�.0��o�TA������ �\�ԝ��I\N�.���nҴ��tc��W���~Wnt�z�/�[�b�NZ���� �*��;����T:�[�V�|�R5�F �88MbO�:�~N����u�S�7v�|t�����L}�DL��7���Z�,�O����L��4�sT5�5��Բp)����J�F ��%��t|n%>�ap���$$���TC���T7Mb��5��:����g� ի����W���/��1��@�0��ׁ����_*���Ə����zZ����1���m�@Rn�KSb�v|��pm�&#�����@*1 S��Ҭ�>Z!RЩT�#Mt�� ug� ��p�h��x�ja�$��L2�N�s� U��x�3�2Kx�೩Ⱥ���w����q�ޭ�͇���>����	�?P�D��^�|�
��!ۦ��L��+�m��G��������篵��D)�$a�H̫N�,^��oN�h^�=:�Nga /���"n /�J�џ|}_^�	@�*Mq��P��OM,|�c�'}C�����̫*��"�W�>5Q𭉄7?C��P�U�����;?7/ՋP�4�������-�t	P�C�
�
�z%T *�p	P��+��m�ħK��N�G�z8�S����.K��:e,�S�8%-�C�B8K54m)�����b��o�x�I^��7.ୟ}�7�x7߼����~ܷρS�\8�/��'�����Cf+���Y�i	@W�n��]�Hk�EIG+�c��2�&)2�mC�ZO0�S��	�Zb��Ʃ#��x^x���D��wT�"�Q����Xb2F��Lף�H�V��ЩG�����\W' ��Y��W��۶�P���nʟc�����6^�G�ڞ�F��+�I�w�p$���̋�$��O%#�!�葩Q��l��R��% �N��3� ����4����B�di>ʟ�d�)I�����c�\r�n+�z�*��T���+�M	D���'#��5���F��Bd�wG�e>���.0iĦ
a�B�&���4��ɹ,��ܣ��d�A$��D���g�P�������28R�L��3����tp�kR��ݗ��#>c	��3|�\J�[�(�J���;M�*��)t$�Jh�{)�qM��� �WJ����VP��$���̶��!A|���(���T?��<�}��iZ丆������w��u:y-x}12j�T������/º"�\�[���;��Xp� �J��	0;I�6H4b�Ö�2d�Ѐ�8�� ���}�UJVOĮUԜ�E�hޒ�������$�2��L�֟�07�b���~���)��mah�:k0	��S�c����'�a�D_��� t1���?�G!t>3G����{�)[���lB��&�
�D�	�6a�;&�����F���a�:��+������	�vp�x�������@�c���~��j!DM���_P��^��?�77��4��T��F�U�gM�9ڀJ���ԏ�4�z�H�)X>k,w�T#Oƚ����'*�Zɠ<�8e�YGi���H�:D;�G�UKgC%RP꙲�TW ꓲ�r6���,�E̅g�Rf	����E/@O"��雲�2��#~1ܸ-��&�����K�;��'-�k����G��X�O��I`Z��:@	I�6�P���1D�I좉N#蔥c�,8'΅]<�K���6�<� ��X1�Ԓ��y7�H���!*-�f��c�2�kOYJ��B�s,��uԌ�4�� j&!B����`	,���& U�kMb�	P��i�_T�sJ�M�V�x�m���q��m'>���*��y�4.h�~�v��12�.z��� =YJ�;�1���y���Dn{�}�1�_{d[�k0�p�mˠCZ�N��)�.����W��>���?�W ��6A� T���������ťW�E�������\���Y���A��#��E7���z�
5W�r���
~��/���'�h���Ra��8��:P鬁����������'?�>���4_>���{�x� �GӰ�"sS1�`ޒ���g^L�� ^4�� ^�	>�3& � :%�O=�k�U�eY���6&������Ǜ�$F݉��ĩ���_oF��Cdj�Q�=��	N�~.=����2 wA�B��&QF�t7���.�����I����e�F��R-\���p�d��s�2O���
�N�m�8�����m�F/ž�M����x�.�<���Cy
����	PO`!���!`*<�ga� 4n9�����cE�Vl.A/��]9��`	?����#Q� �I�Z�$/�F֓�/�K��m�7�8I2ȐT>kR�d5xQ"A����f��.A*��UL��P��z<
�y���Uqj��Dy!.�[�#���o�>ir };�>n��'�P�ԛ䆔Ke4�%@k!��܋�ȽT����i�B(�kmY������H:��ܒ��ɾX�����R��#P��N�w=��� ^"�(i^+MoQ��V���'���-|�-IT#�J,ɠ;ѧ�����[��~�DfA(�P��`P*�RU���B�%>(A�~I��
.��b&�]0���gY��$�R)U��s����sKe8�����X��||�T\d�R�3���p[��1ҿS��8&�T���ϘS��R5��69H�&�&I�9�Ɵ���s;����7Q��n��KH��/����g?�(B5Z��M��4F�h�@��9Q������w:�99���!@s��U����ؾ;�	�ͻ���@ ��G�}Z���&�Q����g¬)f=�֢� �	[���8���	�msqx�l��0e��uSP�f2J��"t���>�#�9�9���A
A�4CC���$?DM�A�doO�B2��j��!�dB��cr?0��S�b#�nJ���UB�����I}���-����a����\:YF�탹ܞAPuho�ӕ���^��I�{1�K��$�Fu��!�6��×���Wo{�����	~�p N��������*�z�S�|Js\��j��q�l��>�@-Ƹ�|�;,�A��	@��. %>�)@ͻ��� ԀO����|C����C��4lj�|��+�P���1�q�H|�ȼ��y*�%�K�(l
@�nI��RPj862���@d��6�x
��n��@�)fld�.]	G�MpH��"$=�*�
.���E���\���빾�	R�؅���݉M��}r��r>�S"�O�B�Jz�/$	P��Z�I`�m�����vq|��)5�-jOt:
@�f1�	�y�K�}���5jM�Z�N�X2���Z��T.��.�;h>-f�s��4�%>͉O����٭�g�c�*|�%�K��/�j^�5}@KL Z���O�}�
�5��f��K�����Ⱥ��8D�4��A��~���H��g�0���-���yz3V�t���02��4o�l�j���c�h4��'�s�~����C�M�U	U�G�Usb�2k\��qj�!"T���)�T��V�>���Qpi�*��4�qt�F?э&��E�{SB7��D��䴶��>����z�{���o[*��bl/���A��@Bt&�u-��E܅�(�u{�U�`G9N�U����^����<���	~��?ş�����_~MP���o��~����������_~�?������/��	^|��֡�v/���"�p&��s��1�x�5�&��5�E���D�=#�NE_^�������4�� @5��i�떊�!R�����j�4��n�,�y��[�f��hx1�<Σ*Ցp�p��P�,�Ǒ��ʧ��2�R/^�uV@��N�z2D��!��}p;z��
�=�e�&��)�I��25��,]wm��T=��ħ3#Kǂ���YFUA	P��:��iK�����ɋ�����{�7x��V�����˟<��{�C������[g�9D�G�؅�US|���A2Q�
L!@礭Ê|l����]8p�*�v4�	���*e&JD4��\�F�>�T4e��m��N���z^�����$.����F��q���*U��Z��F�U@�%ġ
�C��Y�����BhJd}��pl�R�/H��}ۏG�j��1��K�� Mn+b�j*�+����sHn�Dޅ"�],BNG>҉�"%Y�߶f��R1v^+E�B�s]K����b�1	�'�yl6ҤG��#���B���Z3[bL*�286�
'x&��2�k'BZiZSb���J��h4���F�ժ���S0Cƶh �}�Ϝk|�h�L}r)iDi
a�Ҟ�tBT�S	�d9�@�'u�)���9�?��XbNO�gXc��)�)����ݚ��/�dd=�������.($>U3\��I�O�/ =��ס�,Kَ��(�Ж�������ϥ=�Kt�&�(�҄������s1	'����n$����d��S
�*܎�
R���5%#������][��~�Ӛs���)n.î�=(>]���L57�b�\�`��PvB����dT�����E������*��$>#V�>|�BW��9��	�c�ѭspd�l�<7���ӱo�T�];{�Q}���ţ�2{�pd��De�TD�JL�M�C�$/��|N��s_��>��a�j��A*�3!x�`l���@�G����X6F*�y�A���&�a�)Ӳh��@EO��J?�����s�w����1�Czc43jpo<?�Ù�\���n��A�:�:�ΰ!F���E|�}j4�
@�	K;I�'c?���=�@m�&�f,3D� Ԓ����4� �v�'l_x�J� �M�b=��d�(��	2o�g( ����r�QOm�۾�$<�f����s�T?e�[�s� X/��ϯ(�)�4�~>����c-Mo�N���|���IL��x��4��l�8z��8֌���1��Ad2V��T,�&��ȼ�a���d:���BTN�m�4�F^�!4�]��b���9��`ԝ���X��5�I[�����@x���w�*#}<U�3i���)ؕj��sp&?��e蕺.2 E</@����a��Ǐ�[&��mCtJ,��>�6~,"���`Gl�!a�8�8�x�5��%qi��V@jp�4N�Do+F3I�nZ&ςe
�'���D��.����~"�Y�i��y07�rk�� VYa��P5��*�\�ar	���2Ђ�0+� ji�v���mن'b�h�>�>��~���!Be�N5��ai�k4���p�P��S�<@5d�FG�i�!'(xuw�^�4��C�tw�Ӣέί�K_�@m��\V��3~U�5�~>Ө��&r�����h��gMO"е1.
�(�*�eʕ'���i�S����q<�O pJ_P�j��mU��$x�&���A��v�jk���aXS,��3	�Ս)=[��e8z�(�_=�#��P�~k;���'p�j=��=�{�]�����׮�������t�\ĥ{gq�F�.U���(m܍º��n����=���iX��I�R�/vG�M�೩�g2���=C\�"�/��|�b/ޤ*}@�4&Ç�^�����$��V�Wm,<�N�T?=괥��KO�,���xWr[�ښ���?O�Ӄ�}$��O�Ä�Iz�n��U ��.hO����ҭ�Y�}��h�z�O����*8䮄S�
��\����!�P.�_�c�2�f�TنLG���O5^��;x����Û)#�΅{�<�n#�`!��p����	Е����7cuq D!��E�%�)���	?N �ˠ&�X���W���T[��db1�)�>U���i�����$�*�IPKٖ湪���Ƌsm��&ğ̷(���z0/���G�L�T�<n/���.���i�ی��X�VE5�?�����}@X�(�`�:O�Y��	4��yN0���3Y�=��]WJ���~�˟���`/��;
���p<�ؐ�d"%�4!I�H?��m~�~�e�ܖ֢!U�ۚF��Jd]k���4<�ي$�Ԓ�e���0�.�&�\���r_��eb�{D�e���w��^�>�|��U���l5���4N
#�ˤ�2�O&�'��s#�c�i.��; J�����엏u����+�&�X-��~'Q���be4_b.�9E5y�&�zdJ٧����L��� �$)LF7�&���,3����s�w��g�՜�j�2�Ќ;%j��Q2?�I"���O�F4nL@����B�&N�k��r�g�c�i��I�SX��� l۳�{��` ��� �"!�ѝ	��F#�P#P�~jMp�he�"T�XH�.@��y8��=D�����+Ʃ)Z��[4Y�3�!���8�b����>��H�N�B�xO�Ket��'�2R�!�c�uJ����5��:�V�8��.�E��B����I�r�bm�Pm`������<?�#�x`���!6{z����>�D�#�k��{x�����<��M jM|
@u|�L�Q�Qp-�Y�
�����|Z��l�j}^B���+�'��j�LSx��f %>4�j��}���<h,K�Ӓ�
�kCl�O[�g�1v�ĖiLAj�u�l��̓� 4R���G�B�0�����!FmU�h�SW�#m���v��*ҴV�sJ�Z�o���]�;}z�=SV"�9~�B���4�PǤ�uH$V��Æ��!.�c�Dx&��sԶU,�����>-�}<�b%XM�{d�I\�1�Nb�Rɥl?�3�&����& �z���c�yR�$>����e0߹�Y��Z�S�v��������~�]*�z��P��H�N*�F��QL�(њ�vMwX5���-���������:m����u�E>�9g���1
.2�
��_��Dֵj�TF���� *��Ŋq�x��Ը�͋7����ɠD>��ϩx����)�adٟt�y�aD���P�=��G���x����2d�؏���Q������(nك¦��'*��;�}珠��a��Aکb^T�"�.�i�'6�)Nfb./D����S���qY�k�����&/.��y����hq�q��'/V�y���DX��Եq�����ӻ&^�S"�&��R�F/�n"��D��V��W%�M�x<w^ ��������n�#��~���^�=��& -#@wo�+�R�	�D�S�z8��}��篆C��W��C *���Up�Z��٫���v�3�?|Jn������?{��Gԁ<����3z)�� L�����(4� Mۀ�Y���p��G ����Cp��D��УQ�hb��,ְ�G�U}:MCl��4�v�D5��*U��㱌�ahT��a�'�$a�e(/�%aD�$���T�u�T�u�rn8���J�[�H�\��i�ʩ�� �Hs��Q�_���&�\����Px�T��u>Pјۚ����Q�r9*T�Է�P��
�狑DhJ2y\|!�u�F�)��j�Oq
�YH�$�m�T�.I9-!H�3T�^��I�NU����r��#��Ds���'*;r����O�r&M��m��
���d�4�3�#2�/�2J2�)t�iQ��6�'be�]"2񴶌��/I�a�Z6s?��N&�eOȜ��I�I�	s�V����`R۲���/�D�J��Ϸ��K2:��$��=Gd�$������n+TӰ���E>�Yry�/�!�l12Z�y��n�C*Q�ܒ�א�xx��i4?gibCt&��{B�J�8�,��؝*�o?��S�ȩ�G��Dl��m%�߽�@�� h���4�D����YS��@�BV�&x	����� B�B����M3qP�n����ݫ&b׊�)\���D��M�f������"}C��!NJ�F5�c�2�!O(qJ��N�"3���A�f��D�Ts���$wJ_�����c���`�F }^�GC�����	D�!�}a�^ <�����1h�+�|�P[8{�}��� k��{x�������iT���i����$����}a-�ԛ���Z��L ��̕&�>-��sJtZo	��#� D��S�a�\��8C�i�& xZ�����ȴ
� kF��� <%��$:U§�Fǧ̃9vQD�i�P[�86�u���61saC�J���K�"� *�Y�g�J�d�QU͞R�t
@��P�lr�ݾ��+��5��%!ړ���Ǒǳp&�#$�sI�
:�9-�����
�r�M"j��ٰfL�ۧ��&�jꓱg���!6m�S�X�iP�OBRǧ���M�R�o�1O�m�2��q�O�<���1�e�BX
@�|��-���S"�O>-v� :7��*]Kd���i����<�d����'���% �n���Q�<�%�A�i�i��x[�&�gTHW�WSHm��C��{�v�|�nr��*�|�H*�g�̯�4��m+�>+@�DO^�ǋ��Jų���P���~-ɪI�_S��"��L*�ś�}[џ|:Ú�0�d4&4Ea"_�>��M�XJ�j��\�!�}7�;�"�����B,��^��/�6^��m��r^/lN��S)��LoIŨ��w!��gs=��#x��/�s9��}[��K|�0}yq�*�ħ�|��\�0u7 Ըj\	}�F�������}n������Qq���T@+ǻ2B��H`�xL��uh;��\�>��{�P�m�c���lFB��þp�B�C�*8�B��p�������u�l��ҕ(���й��ߏ��&|�m�{���a�E�4_��+ u :�Bf�=lF/�ؤ՘���6bY������b��ϸ"A�'r,
���*�'�"�H8J5�*AUq�JP�8��Y�m�H���³:AkJK,��aD�lG�v����6�e��ŶR���}B�<v0��c��pl�s��M#�nM#�o��ze�� �C/�f��7���$�	��˻Pp�E�J���n�9爸3��"%�/��Z�ZިÉ��("�dꍤ�x�I[~�e�E��q&����-�j;����6u&я}"<O&&ɐ�	,���|�8�=WE֥�p6�&ɑn*��\��u�w��u%Jӹ?C/i
~|�ܧ"�e2��,�\��siK'�S��4��wP� �����{oK��L��I��w�K�  9gIDAT��d-�yOoNE�g��t�NI=��ޞ��4���r~>�s���(Ps�\,RM�/�D>i�]]R��ϱ��K
�v���{����3�]v� �<���󾻑s��m�
V��9�R%XSMW����Ϻ1�'��U������q*{/BY�~��!���uE�JC�E����c�� �8ğ�P��wQw ��S��*�����%@O��a�P�4h	�U�Q�}Nl��c[P����8�~����NA��I(]9A�N�t
�D� t�d���YC�6cR��E��>�'Bc��1�w3�h�?B�ADd�Ծ��_!T�k�"}B'����~XM-�f�D���������R�1��d��e�;&�2a@/L�A�zc3�(H���q���=��m��m;b�{x����n�'��c�HO����D�	<�<�6��W�O��v��~�	����S|a�|�Z�!<	P�����l���6G�z�(XI6��%#��09�k��S|J�
P��"h,�!�g�4��+F�ij�O�S�i��2�}��$�L"����Ʊ����X�<·c�B�B焅Z�Y&ӛ�`*�2MU������
'�I�zd��{��R�=����eh~��
�����Lh:�.�}2Q*P��,\܂��l��t��i/J��d�2m��4�C�<f~��BSbKl�&�9ǆ��qi)�d��G}�4݅ഔ��B�s���8��V�Z���Vd��\�S">-d�!��Y���\
3�Ӳd�v���n�����)h~c�*tn{"2�6�L��}y`�X��Ʊ�~;�7j}�[�He�;��X3�@��>@�4�S��
��m��BY���Eo����s�c��V@��d�[x�y
@U�O��8ܧ �T*�R�|��E������$}y1׷%}x�{��;�UG��KC����B:��O��3�����D�`md}�7�`Jc:�7d`Zm:�V�`Z}2��z*/��4�bg</"��q^���("Sa�=�y�!|���7�\6�����Ln�p6�f�/&}xQ������	P�g?�ۗ��lN�;/\=Pi�k�T��H�'� ����b��b�O���Je�:����/�|*��]�C��VG��J�4׍�Ǳ�n��h ��� �����}�#�qݽ� ��](W;iUPǂ�p�_���"�YӳH�PW�f�2>Aϭ���\\��5|��/��go ����m�\8�/�3���a��N�r}l�j��܄�[�����	@y�}a"��D��f�C�c0���J�	���B$Q�5�5���P5�`5�P�4�c�,�T��|,I#��p�dv��@�.1F��S���a��� 	�Ǣy9��5A�$�(z(��p���*�Tg�)�Te�d��X�=��"�(��{.�BiG!
	�b#�9{x[��8�v#�^>��Wv#�?/�|O���3N�y�"Q�ɤ�)�2��I'8��h�}2Ngi��⹲�³y*m���ϯ����|>���\��D^��ß�����1�p��R���]��k�(�P�b�n祝j��<����ډ�����9s�����\UΛA8f�g:W�ϟ{Y�c���L�i>>�	�l.s���3�(n�s���"���8�Y�O�`��'@�9���s*�P������ϖ2����%�g���������E�	��;��X,�S��w�q��Q��e�<U�׵��c7�c	�[���J��) ����%��I|},�{*�.��)H�%����c/�/�Γ�ȯ/Dfu6�bc�&l.ނ�{x� =���a�4�*�?���xS���hu�"T�����\�o�rl�l�C��@KV��D�c�>�i�� :����� �����C�� R���c�O����|D	�S�`!0����*�Z�G�gYFl.&4@y�oPW#��V�O�m@=0i(�C�N��ü1�7�/�Цi�}��n	{+8�:�������s j:ؐ��ĥ<�<�ް�W>5|������9@�����T?��j=����'6<�z� ��G t�H��6��L�b�������Z?�O�`C�ȴ!0�C��nb\�T�4T=W> ���=@��t�4��M�k(!jO����B��Ep��g�@;��� B\
N�_�T<�����U�s�*`��&<�+w�B�+�+�uH^����ɋ�L�K�>	���]E�n$@��� `v�<��?e>�S�T�S��$@���;b����sUs�NH�V�,MQ�"�����8��2M�2L�b�N|�k��iWd�[��iU��e�a�g�jr+���%c�ϧt�N^�����&�R�ԡ�� @
Mb�G=���i1����Pm�"b���c����O���]���)�ʹ�O��J�O}�!A��'�Y�]z7�)��"T�����j�O�g}��~�� �Aw:�IF��$�k���:��^i�I �]$����  /db��l��A�`ʋ�a��0�)��s�BKF�db$/.�gF���s��ƴgbȹ,������ ���#�R1� ޒ���}���y1<��x1܇�>g���ǔf�2��S�U���)���/Mp}�W	W!�{��1Bc���3���^�����ܫylU|y�ևX�Ë7���.���N��zEo�7��]� zd��gO��K��h/ƍu#B{2.e�n�dwn�}�z���c��y��"�$>��S�
8��|�,b4u)��M�W�,$�ه�_��w��w>~���R<�!�[)]6���>��0(v	ƥ��LtQ�?�m�h��2�!��"����B~\:�<��~P�����Rm�����DrXm���������h��m<�lo����d���Pl;��G�;!*���%��%���OF�l^�'*L�|�a� ��!�b�Mu<�':�㪒��.��)H*O@FU
v5���E��L!J��q����
��9%犰���-g�ev������ww�����M�6e"�Q��2�?Ѭ�<�%�K����J��K���99-��=Cl�g��t.v>{�����s��N��9��0���{���h,��^!�#�[�O@(�'�v�+��ke8v� ^كC�,�],%�vb��=��y�]�V1�G�OfC:��XE|y|_�����Yzn��ζ"���}����[DL֒B���{	��wa��b"�{�����EĴd��"�-��cw�8�W��s��3��s{���y��H��_>Až���m?�Z�b��ֽ�sa?\9�}�a���|�v��cv]���%�x��C��(��8���{P$����߲��-��]Ω�/V��Vv�ރ��d��bǮ ��ـME�! :� \�-@�����'�ס!t�W�6x%!�� ]l��<BtAg5�|��<�7�TUP�4�|�Z1;��%@G�p�h��O�f�}N%k�pd/��9�OP�#�FN�6� e"� "3p�v���v�hQ�uBl�գ��b�����������ܞ���m3����f��+�6�SGj�S�2.3�3QC�:��ta:�9��1�|1��>vp%B{��Ñ��h2}{�QF��qU��!>}�O?b�O/��蹌m?����x,��-ӯ�q[��$,	P����B'Q:���s�f�l7��4���癑�����=R�d�%�%#Mo�ɭT?�'�z&j�>��hMo%���V�9]�ه��k��fv�� �yUl�N|���s1qIp��j�P�(�.'>W���a�&@�Vk$FӬb�q���l~6[��z��XI�����`0� %�m�/}2VĪi,��ȶ�a�} !��!j�(��g�4XGL�M��J�f�����p��������%��x�����*z6l	@{�<y1��=��l�:x}�+`O��H�E/��V�F�՗�2ѓ�^ĥg.A�Gh�F��p%0{�6��������)Q�9�i��3c)1�璺��-*�KY��٧q?(�#�ȶT&McKp��vi�i:߇��KY7�~^�ȹ���OƊ��%2]�y�BX��ً�I�"��d�/gI��e/�o������%6W<N����ܹ
V;W�j�)}>K��v�F�1�e��g3�KY�-%<�������������?���ċPg^�ǉ�ͧD*�2_��*ĀB��Dֻ���� �Lb{���\��;A\�7�Ce(�º�6��S]�Z���2W�a�Z�	Wя{Z��	N�tw�D���8��]���vR��J�U�Z�k�ԛ��X4�RE�����>������?�~ŵ6J5u�'F��Ēa�K���W���K�I�I|�"Ml�����_K
|���SI�lL��I"��>���j�$x��gR�ݖ�y��#b�#:��`�Y飙�!g��l<w.Ù�x5����~=�y��]#�)U�v�@Ƌ���S1� �j��1��L��d��|N^|ާS�ڸ�~/	_�7_�_�o=chvk?�[����������� ��D���'����TAy���%�񾄩���2JUE�x��Gh�'F	%��?bI�>����~o�I���E��A�8$�@�t@��~)w\e�PY�m5T@�Ùuٵ	�\�Q����Г\�7���,\n;�/���X�L�O�d],ǝￍ�>y��o����=�g�G��N\��%p�Z ��E���an��(��A8�܋{U�J��HA��Ķ?�����D��TE!��Ya����y�Ǩ*�"��BxU4P��!|?����X0۹O���V���ߦcaj)�z�0�y6U�Ց�}����8N|�󢛏�D��M�� ���RU�2��_�I�U.#+�U�V��
2�ˉ��)ȨLG~}qV��{����<Y���T���<h(őS{Py�0j;�����������P�zǛ�����Wk�p�Wjq��1hڇç��+Ε��b�y[�y¦�
�
�q$%<au1��@Օj��h@í���V��KU*՗kQ����P�ګ���ހ�kj��R*xn�w��i��jB��j4]�G�:4^�CuG��9���=_�Sךq�f3�O�.�1����hy�N�<�Z>�<���5��Ns��;-h�݌��q���_�FOn?}�5���è��s�n@�5�~�$�_�@�6Կ؈��|>�+Py�5珣�rZn6�j���(N��<s�������S|_j�<�}l���C��6��;��ey��<������'�}�/U��E���Vm_�����������}�	'/5��|?�4r��2�/70�h�ք�M8��`O�~� ��;��'p��(J�������}��={G/�@��z��Jl?�c�9-�T����.A��j�?:�旛Qs����Z�Ԋl4�3�aC�F�w:��_����R~���*����ϔ,��F�6c��	M]����
��W�)�Ⱥ`���Y*�7�PMpe$\��P�gђѪ* �J���f���Y��h��%� �!x��Pi�6���w��Bh�8"t�!��̆��X3�������Y���M�za�5���je��ix*��v}9E5�%>�# %�$�Y���K�����=1lHo����~p��|z�ƻl}]� �}ri�mA(��Kh�����	P³;��9�H���S�ZK� *�4D�ӀO}���S��t⓱�x��q�S J|Zt�S�x~��j���$��qD��5j��q�SM���ɘ��Z��$@:��	���u+���&sr��ܝ�v�T*� U#�N}
@�(|ZG�� Jl�E͂]����3� %����"�˄�NĦT���ĝ �gԷd��Eꐺ����:�2��qC�T�* %8{筁G*K�&8���m��U
��υq"@%22��j����[L<
:���@�
P;!��8�Ecx�Q %>�Jdj %���m�i;��;��c�(t�f��*��Lv��4f�P<��"9�W�4�e�*���Ix�Z�Ӧd�§��MD'�)�ܳ�{�LnDe鴗������4� ��p��P�c�;��d�WS�1<���m9�å�������;�:Ȓ8�{"(��LU"�t�q�P�֏{Z��Lo�ݱ�<�D������Q	�O� ������R�d�N��U8{�]B\:�6��ʶ�S��KT 5L�" U%@�� ԓx8�ƛ�T�$ܼ�L�/�1��4r�D����|�Ln`����*P"����㐳����ٗ˾��GXJ�+�f�Z#4�p��0�g(��s�c���b�i>&ӟ���ss?�L���K�צ�L|6�'�M��4�Dh7����ĥ7��B�F�5�'�S ��Y��\���U������(��Cp
@}:B�[�q݋p�$�d��h(z��	�^���zh �����.�OY������� '�1��e!65���k@]��#g�^��s�r�͛	�3�q�0�~�-���u\{����b\�����E蕰�q���^Qh�rt=�el��� ����G�~��m;��xX�sP�� ��a�C��R���R�A ����i/�����;�DI ��mD�?oxn�����Y��D���" %:73�a������0�,?�����@��4�ԧ �Tқ�՜��UɈ>��c�j=�&I�i<&yͅ(=U�=�˰��>��?J�U��F-j�����Db9j/� �*q�����k��G�;?�}�6���������}�/�	>��[x�;o���^���������5�x����WqCE۾�\���o�&��"n��G���7?{���;o�ƭG7�����go������|���[��x��Cs�\í�o��o�ǃ^�C	���'�|���*�����?ă���o����������������x�y���q/�~w߼�^�+�z	����q����w�u�G����/��;���o}�>�������O?Ʒ��^|�6�>���o^��ׯ�򃋸��y������˸���}�^z�ZJ�y�^��W.��7>~/���t����&^�s��O��{}��Eٖ�p�-������[/s�|.Wx\ο؊��gp�v.�x箵��JZ.���s�;S�Q��s�^�KjP͔�)����*bwuJ*KPp� GQT^�]�x�<u{������{�[����;����)�=��玡�&�K�:w�;�t4��c�!o��mG�ai~��r�%B����ClJ���J5���GL��O�t�f��ބS����h$D�B��6x���V�@Dz?PC�S"Mp�����cѫ��w��q(�q���"}A�<����-iħH$I�����iZ�Qh����c�T_�@f!*���'��V"t�X?�}����\.�!t��)�z�J��Q�3����S	N�猑2_���P��(�7���'������v��ý0� ���GO�z:���v}\`��o'X	D��Mߞ����3jCx��5J���X��Ԋ��2��j&C|~S�Z/y�zl�y"��|�i���\;6�`�$/@��ӉK����iDt�Ө�TC�ql�O�ىO��vvg�m�عp��["�4R��浦���g*aG|�%/�����B����A��f�B��.��H!j�Dh/�z�{P�=W�,e��TEe
��ՀOc�G��(��2�?�L�9q�̅*�B�꥖n ��WT���� �p2�KUŔ�;�R5�T7-��&�]Fx��e�
XI
V¢h,dp!�h�O>K��Ve}� uڷ�}�xy0 �ǂ�C�yh;q�G��T�\��h����I������ ��dJ�*��瓱pU�Hu��4G�*�6_�&��uG����8��i�+�����X�Z�K��uOF�ۣ*.�L$zJ%�q�і
�ĊT%�P�lv���BX:q��@$Kbn�8�5PWBUC.�i��)^��IP*T�@3����Bt2�;��J�2�9�ӼM��uO�2n��p[���%�� U1l�&��TF��#@��>\�#�S�@`d�E��c�؁<n ��/�f�����}�2P��_�����߇8��
.*�O�� �ۦ������g�T9�`�D�)Mveݝ��u�K*�POƻ����*/��2@���I$yI*ܖ}����p�R���czQ�ɋG���@��"ԕ�/C�=��{�t3�J6��) u&@%N�����1s�k�d$�ރ[�}/@�^��,^���X�P�3fz&�	����ы08n9&��YhQ֕� � Mh�EL]���b��@����u#>ٖe _�vF�NFJE��=��]�K?��Q����焌B+ӢD���ح�M/�u	���2�l/��x�L��W�i�&�D,r[rQv��-yH�ME^S2벑\���)H�NGљ�8t�];��W����8p� �>��M��:\~�2��?�F�,^���{mx������{�����!~�����o����_��������}����3u�{����?"�����A�+�5�-B�O��{/��kD��K���{x��G,�K��wy��;�x��W��v�.�nǋ�^Ý�ԽK����:p��jy��9���^�q�y�[x@ �O�~��g��?~�����=~�?������'��>���<�=�������5>���.�"��K�p�ի���U���:_�m�N�>��}��K굼C���������!~��_��O�ꏿ���|�/��u�ƹ��h9���t9*���([+վ�K�8{�Z.6M|��L����|�����:��t^��+|�|.���8|��>�^nRˎ�gԾ�^��w�,_O+��=��f4�V��z����^<�+w�q���*�~�E��Nx��BS�R����X�Q�?��|j���D	
�#�8	9{���;�e��l��ު=8�t�廐{0��iI���MX�K�bY�b�Facj�T��F=����H.O���m�8����a4"��C\�� Fu2�Q"�jej�$$�3��X"Ԭ%f��Q;+�к�e
�z%��6�~j �#��2�aNPU]5%+ƫ�Pi��#T�fI�=D!T��2=KҴH�N���'TU@e`�ў$�v0�v�t��>�< ��bl��:�t)�Djh��`�'!�y�\�_2ǐ�D�t�s&�)�5�3����]2���� E����#<BG텑�#}0z��q���z��>�Ħ�}`���>=`�G�j����(�iK�Kl��Xw����>��Y�<����f }
>m�}"6�UF��~����)�T#�>��@u\���m2Y�;��\��Qs{FjU����Cp�QK}ۉ�t&4�/�i��)Q�R�}�q騐I�ʨ����O�
<�6o���R��*��c/�c	Q�l\(�I��&@=�	���K���. �_�%�m7�ҕ��h�cl��Ϝ�����#��%g)�/!>�2`S������W�N��B�i����k��L���J�Y"�ۂQٶ�]�%Vgw��[����!<mW����,^����Q�OC�S�i�[�[�:�щ|ʲ/$��ѳ<��Y��= �>�2��� �
@�n�ܶ�p��+@�Oh��*�D�mUh���R�4�)(�i�� X�F���F�Y*Q��n"����Y��Jz6ƪ��ng/���nMD(�������x.:5�
8e�wk*��z�On��'���9�6b�l�Z��1��mO�߹t�i'"	�~ĥ�S5�mI%T���:�8[�Z�K3_�Hs߾|l5�
�� T��&ƪ"�LK�VI�N&¯!Aŗ ���&���M�4LYzV�Uĥ S��VG)�*��vU������� B=Pw"��L��uY�#@y��F��sn�����04�uUMq�?�?\ʶv���$s�Js[�=PUO�1{�OY�J�\�1j.��OGbs��/�o��
rO���5��\
��U��$�o@�bx0�V`B���ي�h)�y4Qթ;��}��q0�؋�oB��GCU����Q$A\�}�D�\KU2�Ќ���*�rBK��x&A���[P����{���i��=���!|�C	�p^D�7�!�V��E��q�	�;Ghf��\)�2���F�r�ܨFŕ8~�\���1ԿX����#(9��E(i,A۝6���������~�*�w�q�0���e���DЫ���&�ݺ��.�ҵv��?��s���R���*T�ŉ�#hl�AK;1u�	�o=7Zq��i\�ފD��z�X��ҍ6\��3h�8���\�ڊ+�x��'�&��<�߼}�.�<[��0=������m�s�
��'\���<o�$�Վw/��!^�qo|����-��ɻx��7��W�ʣ{x�[�������u>߳�p��ϑ�c��k/^��7q��mu��;q��e��U�����ɛ������w_�m��*��W�;�Ϟ�G[[��+q��q4��@S�	�5ũ���hP�]�%"��{u��e���>>���Mn��R��u��v���ھC,�R�W}�(���D�J�tԡ��r�7�ǭ�q�(����µ�=
�|OO���sl@cK5j���O�@s��������8H|�*���H��� oo62v�"}g
2�̒4�'F�l*BYE�!<5q����w,Ǻ��ODř�x�C��ۯ���V�W�!�$����%1�]_Kt
6뒑ܐ���4��LWˤ������3�g��L|6��GS�:�/CC�r�:"�J#�r�(�)�PY?�a��T *Mqw������Y��S����
B�	Pi��9g�	�����B�&L��	����Q����B%�|8�/��D��A�2 [&��r�s�B�K�ED�B��(�:�3ޘE���m��ԙ��)(%:M2mDo��N!�&���	#�0�y/������C�y«����	P{�� ����ΰ�UA���d���v|$�|�l�{j=��	Pk��)��� �]�$4�ح�Dl%O�n���vħ������mM�?P|������;iV�-@��>�ɨ�=�m�J��O���|��K���+���V"���}D��R�) �%@�N��ӀOi�+R�t���3�4�%3Mp	E7iv�<=	P�麀ԍ��I`W:Ր��+t���te\r�+�:ei�T}8�4M� �
j�8��y@m	�g�M�"X�,�M� r,�O+B�:���Q�r�)hZ�D�'�Ix���]�����`�$����V��
>K�Þ�t(��>k��h������TDe_w u .�%
��7S��`Qs���Dݤ[�2��t"���iw�|Z���ߓĦ,��98|�O=>'n��=-��c�҃H����"���mg��!�]��b�ʹK�	�T?��5�hM8�y&�ȴҜV��)���t�|>�O���1���'���W�[�N�o��?�0�hT}H�</޷����x�q_;�j���4�t���ud���hy>��9������y2�y�^�4�iT��+�<�8}ei h�F#�J_O��k:��
0�T�hM�-�TLBR�u5(1�)K������ U�o�F��P�^���1w"��H0<K��@�ء"#��޳{�����k3z�w��jZ��up&B�������V�^���܎���װ���o��x��G�y�/į�w�2x���[�j�L�߀�E��'@�cB�z���'@w`�n�e"�'"�@$����k��~Q���SG����O0&�' ��@T��D�VkS��T-QU�L�ZF��T,�]4E3�U�a��k�a&4��d*�xQ��ȋ��<�.DqKJ[w����h|��_m$.��t��޽�+o\D�퓨�X��-Qp<�{������`v �4��;_h�N����G7q��5�~�*�߻��x� l=G��M�fcc�J}u�F����+x����]���u�H0���:^yx�������{D��;�qQ�y�Z��3���{�^�7n��E����������>��~�9��Żx��ߺu��k�e>ރ���;�⣏�ħ���w�}��\�EⳭ��%�����֢��('��Wġc{��p��P�P�c���S���D}�q _�q<�R�u��DKm�9�[;#�Χ:V��D���"J��������;���R���u�[�Ř4Y�4͚�-�_˒��ޟ������%�����ɨ������&������i"sl��M�I�>���,08!��{���
������g��Q��M��7�PоA_'��И\�C���v��qv"��q�-��r�^���	��6���P��g���i`���s�h����'��|��8�_����n���y�ܟ=���`��ﱏ���s[w'z�l�q��9���Ds����L�Za�i���Էա��M]�Q�zU�EycJ�,(�-ByC9NV��E���$T�2�(;g���<���@^:��m�Ό��s�o��
�����=�n:q���rQ�wʝŰ�e�ge_%��U��V���J�iO�j+�j�o? o�~xr�1�p��������"@{�w���6tgmCW�V���
ہ-hݿ���{�ZTT�Hu�}c��W�}IAT�⦮U�f1" -}�����{8�qN�$!�(�#s��0R=���I�޸G������5��rv�;^X���(��T!��I�1�p���z�k�ϒ������'Yb��!���Oy�Wؾ���M/$b�a]<6�_�&�ĳ�b����|gu4��f	[t�Q]�(@�����~����_k���x!��S���- ��HT��f��{9��[W Jt�mLB�&-P��M�jڬa3��O��)�ic^𩏂+ |�o��-
P�ۭ��=k��u�LK�󼪀�;�&醫w��(��_Ox�4/�m "�Ab3s~L��鰖9��,��Zu34�� j���S�74���9xJ�1'��S[g����ȧ�%�1_F��Zܝlwi��5waI r�%D� S������q�ڲ=�%��)�
�|J�\�WC�KS�Q�gl�nľ�}�ʩ�SK��s�܋X��t5�q��"�+w��v��M�,F@���T?%_�6���\��P�D���*tr�Ns���?��٥�M�����e&��:#k	O��Up֥!�茨'8�H�3�a���h�3���i"<C�)�~UO-ڴ��)UP�nk����*���V"tA"[#���l�[	W�2+��(�nJTF�efG͕��d��6���b೓������Ax4`j�I=��l�Ӳ,�Fl�O�~�f�;�2?�X��QAԀ9���܂g���
����q��*�|��ԠCF��>;;=W�\ʘ��F��	OA�|�C�FZ�{�=�g�q�KU!�u�(lh�x�D�)|�T?��8i���4���y %��*p��M�V�&�d^�p�'^ޱ�c� Q�W=��˰R*�L���ʨJ(#�PF0*U�5z��9�Nm�Q��g�]�)m����Qn=!jD��JeS"�d>^�)��ga��@�&��y���)�X1�gS8/Q(%>�2	Pi͝�,tJ�� �T<�|&�	Ę� 4^�c�s�
͈�� %�@���t9��7�:>�3+.s��!�/d1�0���2������U}� � *���o�����o"B���T$d��c�>�w>��gw�^�/�#� M,MG��M,���ғ�c%�� M���O��[�98z� ��b�h.@�5W�� �[�ՙ���:���Gx�{h��?h��X��Y�B���EDfZ�S̶��%�2�㸈�t��ɥv�h��ڏ�3>�P���t_���h�hA�t;����{�������g��Q�lAm{,u�8ZzY�*�@���x'�{�����ȯ�ƙK�fo�s�v?���3ԉ�Q�z�bS��zZ��1�v�������A�������x��O��o�� �'��G�w>�ĽO���Oj�pz14�� 315�1�N*�����>�x����c~���#.�>����c��nߝă��ŧ�4����Rh��nb��k��w���낽����J#���j���Ĥ7?b�6�}s��!��1�sH;9���qܸ�>�s��%Ze��!��z199���QL��G<j�g����*,1�n��o����}T�������v��V8x�v���&�]�*nO'|~;c^۠�<K�)q��
T��}�2�9tt_V���n��5��z}��c��"��y>���u�ٺj��vb�����V�����\=�[�h�
���� �����8��5\V}
��N�-D�%o��[������y,�x��?�|�O}���O�}�*�v������s���:ڄ��Z�#aXqiԊF|�8���h��㿽,8�|��    IEND�B`�PK   �kgU�g<��4 v; /   images/b9728b98-ae2c-4f30-943d-a61b81bf7cce.pngd�w8���6;H��JQ{���gզ�jլ�#	j��R��ݢ��U{��*Jc�ڳ�/�~>����=�������u��}���֠$g&  �w5��  A  � %���fP�-�����
�}?��䠬� T%P����<4z Tm��.�b{ ���]������F�@���[g��}�d�>�z�̰=��h4=���9��ȸ!��$[$�����N���OG�,���F�X(�#�>��_���Y6���3x �Ag�ÑCW�~�t��D�)0W��b�~������ʽ�j�W��h�~�]��gY_/�4/q�;�|lG�?���]o���=�@:}��K���-��?Ϣ��8q=m�r!�(���qc��1k�u�G���m��l5Ƽ�+r٫Q.JR�8��J\�W�M�-X,#,P8I�������ZBjK�&5�5	_��wv�m �6�]AƐ�]0�~���	�.����,6��5,��t�9�h�G�!T��ƃ��*清Z�[߲�RS����{2V����)p��pΘ|-��u�_�r��*W1_dn�x�i��)��gy�׹к���W:lf�Q�<-
}��j���;'��4�*�,��V��O�AG��X��(���|��'$��l������v�g���\�r���QE֦��]&�zi^�Eõ6W� Ћ[�{M�^�&���C#D�M*=`]��Т�;���V��w��l�a'������sq��C��8�C?S-��rAK��)�7V�/�?���dn}�����f�6�%����D�u2;{�@=|܊Z��{���D(���}݄���Y��U���d�T��/�r-�?�.n���0P*��k����5�627��^6������?�"�mJMXH�P�±&���x�&ݠH�^Vh��$nʼ���D��\M�/��)}+S��o��+鹶�\��w��5��LZl�)YQ̱����x���ɌI}���)��)w�Ug�����CG��a���T(�h;krU�F\sޟ���t�o(u��xd��U�% jH����U�Е���i��,/̈́��pn�}!�	���X����E��{j�-��+e^��R�������v_})��p��v7��k�����[����m���zɲ�ɫӆ�/�#��vv�3M��M�8�$x8���*v�
v_]?�5��Xbn�Q�����B]�4�?8�tc{�B��6��f��Ħ֬F�{maG�U*�wY"����љ�PT�-���i�?_o9 g�"SW��_���'g�*�����]���VQ�o�~���Yٞ}�̌�!���yF����>�箳Y���H,������e.�ڞ[V'���{����vG�x�t��ˊm�-��iǶ�a�6����~Tَ��z(J0�2i�)o:��F�V���9�o��1D���e�`�ra���Q�J��j�����;a�<"7)kr습�ZpY����&[I�E>JEE���������f��׆ p����ֽ����Ư�a�96B�ib�!aN���E\"�Ru\���C�m5L�yD�gZ��V��1o�]�[��ՊQ�>{Db�wd���(m���gL�H�u��Ғ熤�eȽ
�n��fؘl�1��b��Z�d]{�v�����zob-6*�;A�A��?�,>�)��	��bg�s��5Z��T�K��X*]�3�`Z:K�a����*��\�X�=q��� ��/&)?D��~!--k�3�49�!�ݍ��������A.��Z�b-�[���?� � _�l���k�$.�o��)�R�v������(<w-����3�Y&��_T��0�>�s�mc.�
C5��E| w��,�a�?�*]�I�ϵ�����\�=���3��#䖔�A�����*��JUQ��r�F���^I	�x�[�D��B��_����~fp�˽!��-d�+]�MZ�vl�6���V|� L��<����7/}�' .B� 
;}-�JG�˥q�0���E�[siQ2!�5k̑�!�8��4<�I`��.�A��%M%ռ�3N��7|�Ќ�Ui��[�+3@tT�H��w�\H����~y��7��W8��rݥ����F��&D#a
l��G�1E	B���O�ɕ��}7�v
�~x�@�Y�nf����s��.�>�T멃h�5��x���uT?�t�Ҷ�`�sU	�Y���e�Ի7���W���O��"�~N��]+�?u�F�ҧO��!cH��~�#����f�8���i��<ny�eb���>
d�M�2C��,�;T$p�`�s:/�I�;kKD�7��}Wi�j?-,M�E�Uyɕ.5(���4�	d枽4��ã�v�{tB2�:L���XH�W�e'|���e��� �t�����=��fI����~�<�Y�]�&bGc��ʯ���z����v�E[
q��|��\-��O�r�P���&�盷����\ͤ4^�kdʞ��gktQU����z?U�W"#���oa�yny���q��mZJ�lߠ�x5F�]��S��95�ʿ-3p�:L�S�F}"�u蝗��SP�����Yy��S����
�S�	JNoc���vGI=i5����)* ~����#�}&�*֕��R��A�����sv��˻�0q�ҁ4�u��C�/��=�Q�?b����A���d؇<�<��Z���W9.������%�����5��0|.��E�?��-�z\Վ� �7R7�(��V�e��?�t�-��K�������97��c��K��f����r��e@�%�rf�`%��C��ĻhJ\�z��#�=uo�&)n)�i��d��K��i����@���j;��o�_$��Ħ�r�-����YM�H�_*9��h��g��A"��#�"�4��r!�|�ש���]_#�+R��wMS{H�$I�r�s8E/I�4L3���I���z�����%"��Ù�Z��Q��j��.�,�!��:�6�͊���̊�
x�!�봬��G�R:���a�@S�ˇ�J�SM��>���5z�BI��Hf����`��)��?������M�Gߛ��O�ȇӅ��q��	��swԉ)��(t��g�s��PQ�O�N6KP�ki[9��WEFJ���R~p��n���l  4���zi�z�
���M�ﺉ^� �;ş�
ȅŌE�RY�%޴��BH�s�ny[DIZ�TN���b�ά#�k)}X�-��l\�$]��4��%��i���Y�$b�0��ȇeT�-\�]C�^����{#Z���2�d P֧�zkT��V��<���K��Y�������+.8�@�ͼ9����S�]�|Y��;s�ɲg5
���-����ɷ �u�����	��r~Q95@�����*�S�6������n
�����\��\�\�e�g"d�Q�gKW9k���N�����|K�#��H��{��S�4�K�9Hx�m���N���� "�Fc�����=��gB�Z�����C�ֺ	����>;.��ʛ̋�.yڛS��f�G�@ڰ�G�uT-EB|7e�.NA��zl���S����7T��_E�^= �`�c�/�h���>6֗��3�֧I�ݹ�<����)�}T��
�Ztg�US���-��_��d	9 t��$�;��ϙ����;-�Y[����t
���Ȭ�4��ʨ��n����4������	,��������$n��T��	��su�gj��T��EW5G�]�8_��ҁ�W)��3
�sl~�.:ʷ���_��6�H�o�������l��s�p���2+�8�}�\	�szlٴ���ږ~��-[�;+\�x��g�cB�0Ʃ;^v7�,�b�1]J5�X0��iTh�G�ӹ�_iJ�����9�QY;T��:�����Pf6�����G�e��)2�؊	C�;��F�+2!�S0��ʢ��? x�hZ�-d��GF���k	��d��2�Eo�P��S�ڧ�����+���.6h��ܜs��]�K]�ȟ�ߗ}?:��n�>�)R%V��Tj�i�i�	/��Īh��IOgJ��^���ĘӚ���
�+�l���{5�r��}��w�ޡN��B�����Ţ��o�#�{";��ɏZ��X���[��wx��H�N�M���E�m�U���P��
+s_�ͻ�<��n�+-O�̘��k���|�k�ǭq���C����uONHZۺj���M��7lKJ�Ք���6GbW$����2�<Ju�Q��X�{5�}u���r��B���L�f�~��Z_H��6spW�®��۔1�Fe���r�w�|�W�ݷ�#B�!<rD��'�=�����c4
�Z�c�]]���IN��^������$L�*o�p�>���f	�7ڡ2W�逭d[� ���,�	��j���kv�T��^-��bB�����({=���ٝ�bIt}�e�ǉ춒J��\n1Tdh�v%;_�
*����_�,�.��B��|�o|*���OM��e�q��j[�rg��.d�-���>��@��BȘc�E�������TˏƮ�:89��'�U_��g��袕���t�6�)N �g�zL/�2�Ç�%w�����~�l�f�u�g�伮�ݎ"��R���A���%e�8z���Id��n��p=�I/�^@�����z��É�/K�=O$���*�4R�bN���!e��YO$�f������Ǣ�F�,�]�۠\��s�h��t#�G\���N5m����tK*P͜������2������-�F`�j�����ʔ���N���ӛ��:Z��cDW?��/y�֚&N��4��Tg�d�)��5|�����l�K�/T�*��%�+}e�xÙ�	��L��%RV~<�9&�Ro�S�܄�s��u�~�9�iZ3}��Q��$�a�C��|��*)�p��bQ<�zѦ8̲��#I��b*�h�IY}��V.x�dPF�MY-ⴎ���r�= �����ȉwT�ӔQ�͍S'�"�Moz�7Ѣ�N. Ց��ꑰ����5�񍃙��,�kʺ���Lh��nJ����e���l�:�<�4BÐ�1�n�Y�eF#l<�H�o����u�KO��4ˡ��Z�����#��Fus��S�ҵ�����N ]mu�l+^�//=����pU���Q�$���m��������U{	����D�����]ை���]Z[qPv�n(�B��V J�Ջ����|U0	����'�ߗ58���'�^��C��N�xt�TI�<�H����k�T`*�^
;/�Xdr�5R����"m����W�\����Ν؀��Ð��!]Dl$�uO���u猍�%��}(TG7�SC�����ğ�s�Q¯�`�C��u G9U{z"��1e��m��_��V>�<�ҟLxM��#�,Ge6�6���M���K�:����W�(oH�qO�i���2�[liv��&���dS$�e��p�M�:"o��VjH���w¥��$8���5O::�B@=l&��ڃ�g�D����Ӥ�`R�l9CE���ێË��_��W'�xO��s�	x���b�ݱ�(JFN��~!v�FJR�S^a8�^4�4�"!8����`U�L�p')q��b�ᤳʜ)�Y�|n�4�,�������J�5������ns(Cs.��q=*ǃ��z��m���t�#�@�1\𐢋fN'�$���m� Y��c�̯/�'/��ӝ��g���'�'vS�V�/rӼ���*+I#��$_����ѥ��I�p4�є��'j�Q1Я�10+h8��p!~'�ô1��P�CKb����0��`���+T'����Kw��_��%v^�kN�ͺ$˯
�]��b�_������T�ik&N�'P��L�� ������ͭf,�Ɯ�9� �ܲ9�)٠(�ðW��0���{��6���dK�(^��-%w�ѽ�`L�

d�.�j�?A�ݹEjif�N7�D���ORo){Pp&�X�4�6���}3Ў���uv�gJ���ejJ��	�(aQ��Hj ���
�y�C��:���,=8�DJCÅ��U�'�1��~���@V��O�����m�R&JRw{B�q��{�1��BԚ�]��FؖO+�k�1zmP6��.���#z�e�Α�Kmz�O|�op�f��É��ˑ"D��@�)���!����q�C�VM9#�����	G��_l�L*8�"/E�'P55�7p���X.A�$�'��3~�VY_�ܲ�
X����!��������w�hg���r��CP]���D��0�����y�?@�t����s��^��ʧk��2iċdl��]^������R�d�3k7gI>�䝒���^�aW���v=/2��e�pT��U����ǉZɀ�U*��߅O:�Z���e@���O�_�K�uRK��ݯb^��ȼO���A$�����V�i;|�ǣ��&��9%�� �`s�B����KM@H옓�n��/h��{�f >B.6M���isw���֮c��ANS$T��0ǉ�/�ϭ��I��/DG�(�P�֑��ԩěW�(��0�F�����K?��T����^����#��KX��TW�ɇ���a�~anW��#A�JǵZ�%j����>'��{��c%Qs�J��(��,i%�w�%�#_}gΕߜkxLx>�'���usʯ`[�0]�XDL2��[&bj�H��{[�e�Ϫ�y���+�W�;�"��
\���N=���!�ܦ!�j����y�q�k9:�(�&��P�O�#\;x�t���euVF�q�ũ�a�!�+������[�;�����~:�q���Aqtc�7��� ���%�U�@��6��:M�aU�`01)�~uEUt��d=U��)���mk�G/�>���J�}���i�muB�h1�z.��\Ԉ�K��<���>�ɬ֑��O_�Y�=��uzP�}��,�����mmF���j�e�l?�{D��x�G�f�\�����bGO���G�G���PM�<C��5L=�# }��_2 �rR���.�g�xvW�(}��t�i-�x%�}lX�l~�4���Ę:���^�8�)X�����r%�PH�J�+߼�!CL�Dڕ!�ݣ\��om��4Qu��:���k2����7G����'��J\���49�&+&S^����HB�"��Q&���.�9n��gr�b�� Už����Gx���\�<�]��<��Htx� ���Z�����[��&f?��>[�N�+OZ��Ba3^i��[���0�f(�>v��Y��n��u��ez͌	��9� u��H��-{�b�(*/];�]);q.� � О�{�ef��ʙ�&Ƭ�-�IALzҼ��xFa�%"q����*"<O�O/t�����`/$%b�p-�����C-�7HܗZZ�����N ��UXAa�BDR�C�5�#L*��X�9 ϥ����>��ح��ȶ ��J�2]�=��9t�f��Z� ��-�����ۓ웲��p矵�f4��uO�\���>����p�13o�\s�ܿ�.�x�O2�x\��N>�Ѻ?������W�U�-�1M�$P��U��i�dt�8�vߋ�l��n�V��T�YyR?�N8��k��MX�+
���yi
��2�F[����Wc�s>�P�F�r��S@���<���Z��ai2%t����S��6��{Q����pd���Wۊ�"c��ԩz=<����h�}K繼���h��l�ǰ�xhUk��6��q��
��Vh-^�bڞ�h��L��0#�AZ �q~�����������Ңh`�U+�x�g�+AOӏO
�8�p\�j� t�(}��e�ms_�s�UF�"-a���Ft2���3��Ha�8�e�+KE��pf���b���a�[�)��!nkdL1��r�b�=�4�}*Բr���(�y�D#!yFy8���D�[�"#z$�����o{����#q�¸�J\�� B���꓊���eїb&J�4C5��L����F�\��6�q�27�@:�\��X�n��t��'5z{H��1>��,f�n\��H���G#��G�Q�qqpt<�ϕ!���N�t��g�S*��~��(��~e"��ݦ�?�����(�E�����%�����Dz�|t�*ޥ�?�+��r�!~�V���Q���d�:��{U�[�>8_�s&���q<�"��8Q��gCN[�u���>�*�9Xa�q]�;���*H=�Dn���`P%J�{u���`�a�OM{���s1si�G͘�-�F}�b�lg���(��z�lWvVC�c��,��m�:�( �I�9u���2}o��'1:n5�^�_�������e�3HJ�2'�X��>_�N�
H��Z�@_��iFb`cԦ��WD�ZG�k(�����S��l�q��~PI&s�I?�u{ �΅^�������T8|5a
�_�(��ȽI�}eD�7�d^���?L3������=�L[�
8XG�[5c�h�	scL�x��AT��D9���¦x�'�9�n��G�Ҳ�7�؍)�o��C��M 1�d���BȦgZ]t����۞~c6����f���G��41�4�%	�{p��KO}�@'-�$�몼�%#�� ��Z!��w�Y�*LN�[�n���YZ-Ci4!���ܾ���>�RΆw͙�¶?
[41*Wi�%���C�r}KG7�grk|�KB��ϴ�4|9����j"yf^,P�6�ƽ��0KJ�8'��p�'�JϾ'3!'J��ߧ�Ε]o*]���e�n�V��62�h��F �GgLC5����(�?�Q�X%���DM ֺ}���ez�%1$c����{)t����<��&.�Ev}ـ��hN>����+��Ϫ+f���4�8�r���)�<S-xH{��l9o���/��"�%�y_1�HI����d%C~$CV�z޼%tJ�����;�t�4^��=��A��2��w�������5�?0tE�Er���#���`7���ۖ�vC5H�����"����15V�KRq��ր�Ǘ���c24L�����n�b� wn2!�;~��-��tVU�%���r��<`*d)�$*�0n��ĵ[�-���8��YF<λRn�"�9ʲ-��1�T���`HV��8)�pl|A�a���#�ҷ*�>[p bt�R;d��aJI
V��q��(!W6ˆQ��jZ +�������kPP�;���P>X������}i����G��+�{\� �E
!X�"�� ��
���}����+�m��{n�>�3M¬^�>�-~>U_��!1�I]�Ȝ��U�N�UYs3E`h9Nd��Q?��c?�������?�+�?Q�E�({��,�l��V2���#Pԟ3�/���h�#���G+^�p����h)�i��޺��&�!3�u���WZ��F$�0�n���u n�7 �{���ӱ'5a^V�N#�{��lj�.���>*�|	A�K��9%}��YJ����嶳�M�rL=P�r`Z��'>պs?�r�N��=;��=0�P���D#���AL*�Iv� ���?���"��H(�f��G}@��JR� �p��i�F�Rٲ��bl^.�ܤ/FtZ:�Qs�b���@�]�5�����!�p��17z�	�e�-�� ��7z�L��X`쫊�ڎR��c���i�O �Ct��?3j�I~�+�s��g�$�٫,��weH�QE��X �o�&M�A
�!/\���l�Rը�#�h�L�0��~p[������ݚ��MEB����4a4'�L�4
A���\S�#M�G��Myg*i�- �d?�ì���fj�6F1��Ó~��<k{�h	Sj?�/�7x�/^�4j
����n!f��/��k�<���9z��C��Q7n�g�������	7��O?��=�����8��H}uמ3ƿ0��}�'g��c��J[�(I�X"����g V�D�&"H�)=�y�-����e�9�י��7�����4��b���,����ԍ#�tX�VVpA��Gd��+_�Ї*n6�8�.��ݧ+H�ds��{��?/>��ݿ>-�n���j	Z#1I�F��c�^�*�9�ȨOm>�r^�#X]�mߋ*ϒ(�l)�������l�"��_�~�A��{`l�Z�v��DD���ө������/�v�>\F����#�Z�}gZ��޷;�D�ڭķ.}�����Wỷ�Iz��1�.|�c!�&�W;;��*��ͪ���<�_d�ޭ��-�R2���e��Q앟R{�w��gƦ�P[A����SΠ���%�ȼ �y�L��tW�(Ls@��ԫ)R��/��{tĂ��Vf� �����ӳx��5�t��9;�[F�>�~� �i'��h`9����M?��DѼ0����F�eJ�u3�<)V�^�������w����b�=��o?b##%{�
OT���bG�i?}/nP���|�X��4j��Y	B����_�v��*��^W�B�*�{���������z�x�]+� �҃���XW����������5���d�eڐ���PD��J�HH����G���x�%�BSޥ �^>�q�������p�Ac�K\j�g��oL*#���n�x-tQw4����Az������n͔Q �������KY
X��)?a�y:�L����|m^�R�{1�}�!u	��'P��d���Ր�;|���{!��HҨ��I����Ã�4�x ���DЛ��^�$��?�8��c�+�S�(Z�}(�M�K��)������-��� ��s�W���]A���b�0�tZ "ԛ;S.;sd�:�����[���]^nj�y*�c�͚���#J�/���.n������d��ksv�o�\P§�ˀC�/��a�$X�-��S"���X���T�b����4���P��<�r�4_ϲ ��כ�gR��'�������'n	ι������epq�D�4��oץY�.]�&C�������$�������vb+�:`6�͉��.���ĨE�2���0H�"C�7�4�`�-�+��\�_��/0�Oo݅��u�f�9���&@ܐ(�L��{�L
ӟ���M>�a9L-�3��q�ۭ���\��v�p��u⎴��)� �E,n��Y(JX+��c���+cFr(ȵ�'��4�km����xɶ�M���E�b[�=;ӭ���z���Yd��yV��[:g���)��e�o@6�:��w+��n�"V��H��� z�iw��b<P����'�x���T
��'=Yv���鈜`b�6'�vm4����'��%�����{@0�����O5Zy�c��8,�{赳;ñN%2d�9��7�Z��Ó���"��@��_E�l_Pv��>�����;y���u�V��+n1���N�H.���/D^�͍tC�$~��=g��YF��X#��X�߬����ѯ��>�D��K;�D�׽�ƇLw��q.�XrV#�6�bNzMn�ݠpf5C.FJg�nw�gwx�GNX@`���2!gx5ك�r��-�9ł=��,�!QF6�NX1IPm(O�{� �BM�=Ǯ������'�G~O��2iNK����߫�_	�H^��-�U��+Ry%�.��)��:ڞ{��7p��a�P$"�Z�u_��!�ՙ?t����:^�Ƃy,���Ɔ�Rl�L;���,W�1M�l����JD�)^#1~K�$�0���<�)ėWav�Ma�����s3���<��[C�N����3��+�^�61�bx��L���?ќ~;���D���r���<p�"<»"�h�к�@
$(w�]���	���'/h:�Q(�D�ƫ�>�q�U�Y|�ᆮ��į�����ˈ+K�N<��Y���}���P+U�:7"���Ob��:c��J{|��H�b��������I�
)�IߑA<�u�\w=�Q���#�/�a�o��n��#��x���v�1�Q��+׿C�R��Q��R�Ə�㥹���(��{��[�دH�P����O�~��C��rc�M9+�pQ��o�t�c/�&��]�f�p����BЊ�MRW�a������/š��bq�-��c�V%���Ս�����4H3о6���a���6*��b��(���2V�g�R�O�f�Yr3֟�~������bv{;����!�G���W���b��#�|�꿌2h+(L�������������������J��M<aݓ��Z�Z��3X����}�pQ>hTG������皿�I���ߒ����%O�_���.У���K�w#��x��/�s�ng��.6��d�Z;����T6A���xF�D���5"i���)�{uW��
+ӵ�6N�I�?�9�j7ݬ��d��+%{��(�6��r�9[pp:��e�SÇM�X>S�G�A�"2҇�������vI	���R�ǫ�e�`�x֛*^Oxo�[�6�m~3O�!��	&�T�Aq"xyI����4/��}�1|ͯcun"�L�������3�))гl"(u@�C/U��^u}̪��|>��������œ~g��C �B�!�J�'���T��!ѹ/H!�ϐ��2�*[�^���n���{|Bś4��\9S���c�a�oQ�J�R��BZW�䞩�v�v���O�c����ϯ5����O��WaWxC.��c���T����;�i���h�M<ȭ��#3���}��"����j�k��O{�:�&mػ<�I�׃�m����}E�W��(4�9�p��U�C��g�PaO��-o��Uc*��pJ>�|�kEOJ�N�[]��M<�'!TH0�o����l�9U�P��M�hX�{�f��JM�1jw�A�(���14������yg=y3�9�mB���?���- z�t�r�[�8;�3:��M�����rjZ�c`*��C
`L0!)(V��&��w�{_�Ϸ��fA����l�
e�~�ĊIf�P����K{���`�T���x�2��5d�r>����y|�Q����֨>Ɲ���Ȯ���c�/!C~�c�m�#�IC��>MҁU�A:��c��a.�FX07
�";�z�(��6�t 2��r�uu��l�h$��,Nhn_�%'̫�ɍ4\�Y1μL*݆����vH���@�nVI�0���Hf����8M7��K��,z�3���Y�=�ދQ�N���^���@C��g�������|�A� n[�*�]��B�=`1
��k(���Q�|2Il@+UG+�-Ƽ��E�A�!�m�X�@��V��1E�Ŧj@��M���ɲ�D�>$��"����*b@8B8U���d���z,����Vrc�w&����E�,pr�P� �M|��}�w�@�W!���{?y� ���Aˎ`ȵ|�s'�W�-���ŋ^��&bB&��&vL=�Fu��w�Kג�;�d����8�[�ݦ��yތ����l�d�ЍZ�� �S����[!�N�X�6�w8?�gQ=| ����e�R���k�&�~
�x1N�sZ�<��E�������C��L��A�)&C�@p�n�e9L����s�=��S����P=�Yո�ԣ�Zλ6=�v۳�z���C���%�2Nvf�f� �2c�)�m�8�BE1��.���ڙ2%�����%1b( o!�/�l�Fq0�V��d1��V��o��zWDF�"�]a����Ԡ��jx�Չ�xt2�_��������c	�����9��������hxE�6�X�Xנ�*�A�!&��:��zZo���2!6`3�F�	L�S.b�4�ר3B����!%�-9N	_&�ş����(h���N쾯��}��/b�ܤ>%��u��Q&�E�y������Q����MU3�t�atT
Qz�H�	W��ث��?�i�����z"��� �2�ƕD+����T�ֈ�BJ��q ���Tf2G*��%��VW�ޓ��|�L��jH�P�Vy\j3���w=��`N}i�A��PSJh�?�{؛"1�BԪl�kQ"�>�ǵ���~�l�k!�^��S�k8�N׉��Ҵ��r=��Q*����*�i�4lw<[�.R��#�{!���*dw/��%�?I�g�n��)Z/�$S���X�y��KU9{�^6�{y��
�8��9�Aa$ b��xF2\3e�Nc��I�yG��!Y|��"Y�;E�}{<_��{�[�Q5��	�K����&��|g���6�Gd�����(`�_���z�[e�p��;���xt��
<!:弰o��|���}�%k9>]��V�zz��{^bm��,��Z<eo��,}�$���䮛�0.`UJ�A[��֣7�۪qbK3��Ը-�
1�� ��#N*½�zU^�n��Zir�ߢ�����G��Ŭ��֭u����URՈ�5<#��4��+�����c3�$�J()���ŧ�)�P�(��\���Uj��0�����*�n���Q��*']�����Y�In�[6���0�|����F�l=@� ��9Ժ����[��""������py}���:�;��V���Τ��?>��TE+����|�jA�i�Q������kM�[��iڍU��d}2��R�C�UK1ￛt=�%��X�n>`N}��u���M�ov.� ����E۷�CM(�$Lsn��󊓏���6(�|����,�����b�ݼ�~�����U�/��gSL*���H!BMc0�ry��!Yտ<�|�eȤfu���]��$":�IvD*X�^���Dt��I��ơ�Pl�P����@�J54��Ǖ~��e:����¥�4���Yl��jT�:ȅݤ˚�/������[�*��h��uս��{w�Ѿ�1��7`AL�g\�����%��d 0�L�/���D]5�;�\Fc������q9j®���!�a���`�C;��x�㣢~�G�K $t�IEn�WQ�
��pp��y����E�Q��x�\��-�	��U}��PF��D��0J�|�<��m3��R��(H,�������a8����g�e��߀$e�Сga���q�LSGoc/� PU�f��9�i��P��+��ӕh�㡞Q�4f��0"�S��4oR��G��F2�B<���`v1ӛy�(�[�94FȐ��W���*
����D�H�<i5rz��� *7GQ��u�G:.�?��I����U�4�F͟hz��o���.��;�:��6��O�-��5B�M�(r��J#�Y	�ƪl
q¼�7��A����V�����a�!�y�	���wj����=O&m�4&h^kݏ�s�mks��-o�t�mo�nb��[L���:_��;0j'*�ۺ�b�!�9%��1�>�|F?" w�K���δ6�ᱺ���)W�en̢�}e�cJ��c?-)2��s
�D"K��)�������*ΖiKn������i�U�������+�Z������'��r����^�=��azqQ痴(�;�㖇��L��i�.W5�����ߵ���Q�� 5M���p�/|V8��Ã!�#|e���'S�����Ra�æ����u�d�v]��b�L�4�,�����-�п�-'0��t��~Ar���`t�_�?��G�g
���;��_Cb��l5�� C�?���ߙj�4�����ws,���X�`�zT�]VSb���t�ڼ_�6Īu���p��A���Kاp��.�oaS��<��K锤��R-��Z��k�,�{�����Eu��x��r�q��M�Vⶤ�ϗ˄C��A=;Y���	Iէd�D�D[�]ay�������q+Ye����p'�s������*�B���Q���>�U���dR&�mf�4rI�%^�[�����W��?�B5�X�h]���d*r*����B~��SG�F.A|^ڒڬ�*��HH"e��\ ���1c���FP �D�~c�Ɖ-��y��~�:n�{剈�<�ڣ��RR����)C�$��!|�y����&�8� �P�6ܦ�R0 L�N!���X+r"UstX7k�q�E�GW-dڸ8x��h#O�p`N|�tקw�$����Fv�ؒ��$01���rS�O��i�C��|�2��B��Q0�HnȮ,1�MO�ƙ��yB%�*&��G�Taߵ����w٩yHV�p�$�O E��^j2U�'�ye�w]`2�wb�uRߛ��6��Y���lf�b���`� {�&��%���xFM�2��3 �U�&'}$��'�C*���҆
k_� ���cl�u�a��6��)�p���K��?k�9-L��n�*^���`V_�{`����}���9M�V���D�nȄ��s�nh��I��+*�Xk%J.�b����M�k���AV�/u	��yŦ·���tM��u/�b�%���dX�>=1��H��-�]��_<�M���^�ΉѝY��W�K,�)pF~ *�9�7U��̢��/qʝ++���\��)�2r�p�����[���{e'cƸ��w���c�(0Bɚ���­o�����D������������M�l�ם��Z,I�>��.��.��2��7��a*pu3�7	�w��ٓ��L��7\o����3���щ��F�%Q�FI��E�C�Q��-I���	"j�B�N�����]�8k������y�}�S1_K��푏@�E�ty\C����m�4F�mA��ԣ�9Y��A��9y0�Hof��2>�)<���@H˼j��r8��V�1?�X�Gd���k���l�M��o��љ��������Y�Vo"mK�U���mq�@$�pК��c7��K�+q�w{�7�õ�~�NWp��UF�6aw,+�/B&"ٟ�V��q���c?R��P��T�	g�/|���J��&I@���Ɗ�0�){��5Rƅ��d��RG�A4a��cp��T����>�P$݌��F
c��$x�?����O��������3�u�bá 6����*V!�����wvY�l�uƂR�Z��<�P{���f��`�B�3ofU�0{�ɧu�fS�le"y��[�J���z�2�Ǉ|:�U���I�nRb�W��d�?a��x{���0����~�C��QQ�Fx��olR�}j^m���fg�0�ד��6��SKg�s("G\U[�*E��ѵ��ΆQ�ӯg�st���R�z��1�*�?�,�%�J;�h����	��aE�����ɛU;�0�Q^��;���U�nL�q4P��ƥ�*�D
R=1w���q��'����ڈ n%�
�R�������i	QT�����H ���G<p~�ي���s�0$*e��T��k8���)�{ ����>�MD����6����L���;��Ǘ��S��;.�� �F�G�����hl�2o��/��?�H����Q4�������<�}s�42�n���g��4�PP���ޖx��A}���p@`[s�Q�a�L���V]�*3�zρw�b��^^U�(es�X�d���5����V��B�C�/*��y�eS��ԟ�*�����IΧ��b.�Q(o��V}w�0n6!�7�S��t�*n�קj^��G�ߔDp�Z�C��m4����9]}��R��u�����ڣ� v�n"�d�'E�n1Ou�M'Hq�,�Ax���K_]"�J����e:0	/��I���b"�������J(�˗Trξ��(�M����w�\��LT�|���@"QkQD�XY��y������oE��:��g��t�
��S��^�{��*�:0�_O�{���X�h	w���m	��-N���S#�c��Ŏ�9�O�{�=q�ho�2���5��\1!�|��ź!��#�8��vգB�agB=���(9��Y�zۺ�|�TP��_���-kDY�Mj�I���\�:HO^����؈A�0��C#�}cs�¯��U���#1	��ִ�<#�a�xqD&*bB�4���sOHUz�<�c�ÄRS�����]���-�7PW=�-� 9/}u|U���|oA) ���^��ȵ�y�y5��5K��(�,?�#Ǩ��#hݞoOD5�`���6�w��������`o)������u�w~�����׏�h惃D�fT�G߇�u�(q�SGb;����#QC�2;���`=}/7Z����(��X�����
&��C������-)9�#C��n�y����",�/�}
_�_�`�A巟Uy-oo�:�a��9���Wr���w�NX�gl�.^�#F��̣�u�p�c�/q`��߅����Se�y:�Fp��,�gUy������f;J�B��kp@9{��xnG�EM�_8�{�!�\��
�b�aߖya��(�[*	r@�@$E������ta��1�/6	��u�����jtΡ́W3i_ͅ�:0��{~\ôW���waT�A툋3U6�8���R��L���D��3b ����){�ƕ5Ϭ��VB�Y�?~kP[�8/6D�os��$�d�AU��mG^�����F��t}�p��"�����px�Y6�I��Z��t\�8~Q�����c6ϣ�����`k�H��������נ��i]�^����<�}�F�J$2�)��[��b�`�Y˷�=ʑ�*H���U^�,�=z�á;�Z/����)Pr\�8u�	I��G!�u�
�b&�9��^*�����G���pmwٶ��>Æ#v��·3 6�jq�vd�;�����vÑ�}�{V>���.k��aa�S*���~{�{����
N�0	-�woH������u	�Rx1/���Ǫ-�i���(k4�l����������������*~̢�������7�WR��~��A���D`OC|�4�$N���T^U��6#"զ7,�8k����-�(�ok�~��0i��Q�Y�W_v�Ϙ�i]���˭9*�+�1F��Bc��&��2MB�����`O��#��;��D�wn�S��񼋸 �����̧��y�!�@�Ǎ^
�ќ��G0���kn	��7՜w����t*j������^2��~����ܱ�{9^��������=FK�o�ʘ�D����-Cם�LI���V��<�^vl���&��/`�F�\s\���2&����ڭ��3�(��^�����=6R{ɽ[j�zپ8?���xW�z΁*9cs7��5���m�&3GKA`z����M�O(����*y�K/V�i��A&�T��g�-uV+�t�y�C�5��
r�j,�M S�D*(�N���7}A��!���� U���V+\Io���c6�XV&߈����za�,n�t�J%��k|>�E����Sf���at�dH��z1xD���2B�KM`��p�0�k�PʍW�;�w�su(��f���o��O�Y13��G�1�7?"Hf��VڹML���ՒA�?��cI������W���7�����
���d5ዄ��)�� �9���So�g$�|^��^@�@cj=��X��1L'g!��`}6����!_�x~!���[<��}��L���7h�\����S��AB�id�
�;]�C�x ��Ja�F��I�86N�@� ��(�se�+as֌�����K��|�2���c8z�t�s&\�xv�UUAu�������2��)|�4��T��_IPT�r���NU�p 1�	�a�X�B5�1)��ww�q�Q�>Yr����G���� �l�?��b�����?jjV��]�ãu��`MH��<�n� �>���w���aD#h9��1�N��TTwy�/! +X�_��b%-�o^)���?��^�汹Ɩ�h*�����9����<�6!ז}yM�����.�oo��u�Ǫ�)��@; �(5���=�H �U8�m�Y��"ȗmI��>[�,Ԟi~Ȉ_8$�C��9�Ю�P��R�����#���3�a6t'$M�jn���ފ��v�t�-����L��F ON�K��AUq�>�O:�H�$gY4S����_c�=!���/w�W�h�&+���`n����j5p��j<m�>;�y{���N��#wY�j^ք�K��(:��~٣�Y34Ca��Q��늩Nv�zn�Rkp�u�v�v�RK�Ą���֐kF!+���O����%���C��SeH��7ߍϱcF�Э�أ��)�U6A��cH��U�P�R�m�;*N�������Jzz�'����2��}u�nK�)Ҳ���ɘ���;�v�q�,��ܝ�C�����ÚQ'_.<�}� ��P�w��\��&�v�r\��"�<�b� w~��R����ZA����m�+:UoZI� Oj5Rd UU��+�V	�?rm�Щ����~SϾ���^!�ʥ�E��1Ռ�Jl����(�U��_β"�[��"e�7�G�;d���
��έ����c�Z��B�j��u���צ�~B��]
x�^����Gfu�1�	�ߣ�o3�����	�N�5��t��onV��X�8G�5�}w��'o메�E���{5}p�b�*ؗVv~��v|�jx.��6�<1��l�����п(�|���.]��|3���ws�.l�ܤ�S���[Re�C��}����,m�C�&���v$x����H��'�,��MS���<�d�OWw�݆���t6}� ���X�\8��ŃS���	������b˹̢jS�łS[ ����J�R�������V��W4k}�	q�%\H`��)4G����|��|���WM�k/���c����c��,s�F���.�r��h�YBD�.�a.,�����A�Y�\��\bSs������,�?�7Ր6�=X����y�^u�1/���C������Z���Ib@�oe�-���:I�r��_i��q���)"2Ÿ��i�U���$v�P��Y�[b���H��}�x1II*�&��n�S�R�ֱ���4��g�=S�K�����8m���������<
~7�
��O�B��e<���~,�c��	$������xA,�t�gZ����/�tcn9C�	^��˽?w%�6�#�������B�&��ЖdW�o�</t��vc'�m�༔�ƫ�\:���&[^�o�?F\
�bB�� `��ҎK]hڏP
8�DC�\޷?-�N$����>��dvHl��kr7=��B�1�����3X�x8v	L"��+��@d��`õ���,u�V�}�tN�mX�C����ܟ)L��o���/����2�LF����o�q��e p��(��;4�qr�.wg��Z������� �V���+��O��o��B=B+;zZ�G�=7����{��ˀZF��ym$�τ��X�mS7T���2ɲANv|DF,�1�2���"]+,����
e5u�Ӎ/�-o��g�D�%���ʹ��\^��wi��R�B��X>w*�B�Iݕ����C��F���W�Y�˶{`>�0r	�յ_�ؘ�no{{���sl
�>���{W���b7���?<�����ĉ�u�vS���q�-��f�D����F�+�4L���lG�f�����/�L[d�O61nm-4/��ذ���a8��t���U'7"F	9�$f
�^���6� W�t����5TtkW+�s�L���p-H'�9v}ID�E�	�*C�o��pۢQF�y.���)�?|�!�����P��J! ��xT��z�����Z������U����/�?3^�4W�}�?�S}�ʄ�:3ry�w�y�|S"A���.�b.#���le��x�ɕ�H�.HI��	D�&lt�7XԄ���.��xȅ�Y��exZ�b��,���JM�)�4�r�M=�p�L�> nA��
�~���y��h4�>՝I��q{��X|�	ז�/C�0�u�U��,Ħ���} ��;�=89e����+��)<�yE~xsm���6:Hj�媆C_�{4�`����z��������H����஬�hS����_��lk�K7ZjNŲ�̋��D�7����k9����x\ؘagY���\���8n���"�}�Dn`Wq�* ������}M�x���K��I@ئ٢���Q���b蔚�j�R����9>�^n2�����={}?~�(yL��僮�<67�.����X�6q�_�q^�p�pl��.�ʗ`]�	���5��d�>F��Q�S��=�(����}] Pxݘ�^�����zp���v��=����\"��yM�#��972{��Aw�L��M��x�.�j��g|U���|�h4}ۙk<D�X���q�&�W�X�<� �V�2�'���3(y����jG�m�ܟ�__�$���o*��Zҫ���J��5�p�F{�ĴM� �`�ĸ�T������a�*��` �$�T�}uaN�5ċ�o?W��(��`i�=H��a!nt$վ��l�{�Ȫ�d����́��Xv$O*®���;S,7������V�Ȃ	ë�{}�#�qm3�N�Se�.�S1
ۈE���f;~����q�0�N���D��>}o����$��m�&�d6
���u�� ����w�`��DJ4!����im�4�(��>��U���ݞ�uj>�5h�R�bپ�I���~�a�e���J�-%���GŇ �'�1���%�^Wd���y/2�I8`�����8��N�-v�4m���~g��Y�ǏMwҿox�[�u�W{���w<7�q�H��z9�@�/����R��ҡ���u�����3��o�)�@�zv���z��'}`rUߟW$@y54N��yF���p@@:1'bU��ˇ�Ŧ0�@��ޗ[|-ވ�f��J/	�#B3�"����Q�.-��!��`Z�WG�!ٝ�x���X��1;��K�n���zU�/� Վ$M�g�L�� ����v���Ľ�q���pZ����M	�v׻I �[\�Ե�2����7h��6
�����65�Mk�DN�M���������Ş��3�3S-�1ܻǣ��=�.O�,:���%/`�P�	����X6i��a�	ފ�����g1Q�XɬE$Υm#E��m����5̸�]��`��W�/�����Y�+��
�.����<lF=���P(��0�%+��Va��L��� 0[(7	ܪ��LnVx�a�{�5'Oy%|1���DC���5#�G�y�_��_RE7�"%ܳ0^R)�K�?���\�V������J�f�����3i�u�N��e�R}��)#���C"N�Wk���#&*jX%ܟ��\ϕ�0hy���V=��^�r˨�zy�����! q��_)~�൭�����W'A%�nnop��Bu����l����ꀳ��ڦ�T=��|���cEw�@��qO�k"���C����y�W��C 1b�mE�?�@���h�[�BO��^�������iI�P�R�)J0N+[F"|�Ku��Kم<�����OҗI�uH9��~s�ON�Ӂz��^W��96�FFǱg{��3�>����B�h&Fr�=j���>r����!Ow	�S�N�'��M^�v_��j��x3{&��v��f7�����[�e_j�}��Z=X!�AipIs��6k+F�p1(�M0��7@�Wl!�q�g�z��ڸ��*��T�^HN�Z%ו`�Xï�H���$Mdf��������\Xĺ��(jSsw�����[ ��ִNU�^�F��&*"3FQ�2(��C�8�Ӧq�d�]+� [���ߍױ6=+���������7�c���,�D���=��ɲ٧(p�l�๳]R��].�(�i;ixF]8C��va������ %ad�l�d��e
����@2�鈪~[�S#��z���i7����:�&�c����[U�MU4���;����[�o0�jE�y�%ɔ�Ҹ}��7s�~&�^B'O!ɮ��漰PL�#�������3wy�e�T��kj~3�.�Pm��#ˈ!H/�%����2y�a]2������o%���Q�������7���o=
J¬��6ܟ��T�H�2o���fG1��ۜK��͈*�<�~w���b&',Qfʆ_.=0����8��O�?�--�M�	��}j�6>�*Y��\�Z�N�l����Ǒ��G<��<���J��dZ�����oU����KKj�K�ߙi"z>��g{�L��\����c�ĩ�(^S�IJ�NFY<����#�qS\��卒5rn��p$�Ɓ$�������8�-�]���K����h��}n�6k�.���O>E��+��W�mN������/'mK�� ��v}];h\��fpW���L.;������k &���e�����׌PRv��l���P���r�s�k+�G�"���L�q��s9�w��<��_�&���i��*
��)��W�d��\FF��F8�$L/TD���+$��kv8?�Ja�s��B�C�4���6PƂPbQ�ZY���7I��Ú�r�xA�O<��BLH��)W��)9Rɔ�4>����P����r����/w��Ȋ���j 
�b��i%p��'�M3Y=)5����8��f�'ϕ�����X��D��������ȴ,�h�3<����x�@
���wb�@c���������}*�֠�T�gOUf+hg��xs�̝�ck�.�w�|�F��C��e�������>tZqc_������B�hpyz��KJ���+�vZ�vIb��J���e������ri�&�����'s�/���Foѝ�`'�:Sc�W��:���GF���QFU��uǗ�2A�_�<��<���m�����l���Ԏ'���FA�n;������#�?�ɤ�]�F��8y�Vk����$bK�H�J��C<��N%։��;�[e�;��:fZDʵC��W���R�z��od*!�4��Q��<�.�/�!9k���Y�]%Oψ0��{NJ���LM����gp�&j0a����1y�ۍ[#a�|E�����n��K�Td�8�i�Fwr�'̰Wx�d>����GM,ɧ�ú	+�ixB���W~+��O�}�����K�!�1~y{��"ek�P9��G^�.��oJ4ΎBX�9��$��*�9/GTw�8��k����Bm9ݚ�>A��L����LR�,s�jl��xTL��L��^��1�>�>Gѱȶ�|�����+�a��G_�y�_��~�r��Θ�5V�77`8}Z�
q?�m���Q���@�%;4�)��L0�;��U��6��Bw��Cv9ã�Ϗ+��e�Y�����75�V���m;\r�э��{
�|,�j�C��8�^n���3
�������k�I*�$aV{|Mn�f���>*@��k3�O�����"ԟ^}:�#;��%���z��R v��[�`hV2���-B�D:@�Dr��˧a�9�b��
�iL!G m�p�4���K��3-�r8[9�3����ɾ����F���O�?U{G:���:xg���%�F��-?����O:_=cnzX)S�z�MC�-05����D��bl&M�ب�H�׋9��a�p�NL�7i؜w�܊r1��Rsbp����8U��y����6�N����`!FI�b;9�*����xª���������?9��@!�S<��u��:�T�E���Zs��M�p���u�!Xf�r}b'Ǯ˨ѷ���v~G���&�c����D���0�L��3[�Nx3	닥��U��U�EtΨt��a�7�R�;���n���o�3��%����}0��>���f���~M��?����,м]|�1cl�zs�gz����ڌG�ړǼ��^�!�~ÊԬ�g���o+qh��&���tZ��z�Yݫ�k<o�(M� ����$e�{�_T��d�:�M�<M�6W�j�x=9m�z�H�3������#ULE��������U��J�t�S����H�d�	��0��e�3�AQ�y�H7B�s��8����`zkَ��4K?3_
�@?��83{�,��Z|���6�*�[���]jŘ&�L9z�F?V���v�a��^K�A��.�u�ܳ����y������J�Z���<�Y��!����@��'����"��]�	0r�� 0SC.����:>�����J4���*�H�	��Ü/���.����^�άgTk��>�0��ﰢѾs͑}N[ࡧ�
�c�c,����o��myX{)Pa����Z��o|�=U�����Fߘ�c�!�@l��ʁm�J<y��O7PuBZ�^�$�&�0���RS�;~�5�JƏl�! �[���6�>}q�w��|�" 	y/*x�'�c�U�ك������?K�"W���w�+
(�܈����s�����bG	��v���0��<�Yh1���WR7����Le��z�EN�tZ�s�8~Ϣ��9J!WgT����[^	�m����R������٪��`G�6�`;PԽ=��]uJ�@���1�K����:I�r�>�M|�������y�A��������/��'��Z���0�@��4�ЄTmWV������W��4Q؄O� ��э�Ґv���α	�w�T�s�v��>*1��x������McѮ��$��G�^H�FQ�҂�ŕF��8�QY/ui�Բ����k�)�>���r{o�[�D����z�+땷�,�r�� 0�c{Zf�2�;�V�c���2&r��TR~��Q�Cc�װ�� ����PH�e5�7LX�r͕���s7: 8�~C^�C_��&��37g裡��~�0������fp�K��v��*�g�V���[(����E~ g@�Ty��a$���=�N��Ҍ!��@2j�bu,�������=��a�!�HV]�.�G��-*���Z��o$�O[��;y��׉7@���S���̰ϫ��և �텚E��D�V�?�nI�z��楶0�<��Ф3pW��ۀҳC����j���A�Z�NW��Ŏ�E{H^�w�$���Z���7E����{&�N��7��I�27�bz��l��T�{�u:4���B��-')����V+FY��Y)^��; ĩ�<���� ��p���kO�5*����/����UW������A�D'{��hda�#�*u��_]�_u�x܂i�*�o]B�*|-*�L��.<"�`8(�c��@���l�:����9Fd���Q���՞�J���AП���i�� �V])R�V����1Jp�4V�%lU;T�k��mP�������4��8��� �y�ɜt���au�Gj-��L�wg�c�h��4Q�.�-�Vr��l3����p쪪�x�
 E�I�R�P�akz�-����"�,��FVD
E�tN/o�} �3��~���&x$��������H�R.��sEw��7@�5�k!{%���>�y/���p�y�6�t �4'i�r�˓�b��O�����xv��'�$,�n!��w+�&d_vN�ug^H�Po��P��,�-��������[��=�&4$S[o�E��d�R��`j��Ȓx7�ތ*����&��gh.7:�w�Ǣo�lK��7���(��A�����zFz�R���tBd�������;��f)�ك��̴����]�Lx�힛�"蓼�
?�� R�Y֫���2��ʇ-ur����0AE\b�尹�R&�};�z���e�n�'/�ǚ�?o�����l-���'b2b�l�6JW�zF+���� f֧h�c�s��ڴ^`<���[�hT�vdsp�ރ&P��&���o~���9/���B3��@qd�>
ۚ��EAN��@ř-	�_�q/��/)�{�b�;ad쨨Z������d���J������Y^�\$/t/�֖�dd"lܟS���TW���<y]?��G���+w&�����r��FCG��H���o����n��Z�i�Ɏ|3a��4<ݚ
�
+|�;}�a��1����:7/��4,$�>�#Q��kB�(��GC�N����	/�A��p��-��t&B�Zo�l����,�xZ`����^��9��[z@�L��>�;�Ӗ=��L{�eg���g��=O�~��<Jd1*�;TR��êT.���M�xz��/�Fxl�!9��'��RC>Q�n|���~��Ha�a�Qfp�[_�娴濳���v�n�D}��\��˫gZ}ؕ{����uI=�j^|ȫ���������p�(���Z������g:��X�� �����â`R�ղNS��w���b�b�7�C�7*(���M�n[�d����?;_�Hc��&���G���|
N��_�x]��~�ǁ��R��wp����(+��Ȧ�ቲ�C�}�K�Vn웧w)�M Ҡ�
�� N�.)|�M����.��2�e�zlS8y�	L��6��пL�y��^e�W�:�֣oĘ$;HL�t�.�惱�E-F6���G�y�^��&i�?������B�^� T��/.��Rt5�n�1f�ҿ'L��"�D�/?0E�e+�B>���g����>?r�p1(qИT��f�2P�"b�*_s,K�H$�Ѿw4�J�X�,��y�{�FsR��TIX-֔���|�&�Q��	���Y��|����B��*-iUi�+�,��ۺ
�A޾�����"�p?���/��B�����NJV�`�
w��3�ų\�gӅ�*�3���n�u�K�,����c2���"I���[��a�ʢo�^+N��@��6�4w�>F��=VҊ�jQ��f@�sqХ �D����x��>�6��АR�j	�-8�r�I��QtQ�*G��X-�l)���ϑ�*|�����c��t$vS;<#��]��5���T4������1�u�=1�dJD��e����V�b�5c�m�����焄�e6��t?�B�fw��&��3Wl�[d�a�ԇ�n���WhY;	�<-U�'�gLO�We��`����]��Sq8i��V&�i�f�$}]���K'?�9�P��B�H3kj��������\���Q����E�&��%��ˇcz��@5��������Z�ܚ��yB=�;����� ��ת�I?"�(�?t��_�����}S}<h��������xT{���I��E�v�R$S��:f��9��_R(����o���;{$q���g�|�0v�c�؇������u�N��D�t��}	�n!w�;݊�(fL2�eŋ1�Πy��"P&z�Q#��:�޿��m�G�e�V�`���%@�5rh��(x6���Y�D��dm���Ly*=PU��a��v��M��#%�������ͣ��aGJItx��U�w��)���|N��������*ږJ�ɬa��y`->v�#��a��T�}y�tϳ=
o 	�C�<�(k��w%�y'��m3��̩~�0�HV�m������)��{��h��G{E�qR��/�Y��}�s���4�in۝5^I�=�����n��tm�@Eh�@Xu�V�Q 5Z���{F�?�^���z��e��߫��p\v�
0P�'����:g� ��A5dG�BҦ ���7~�> 0��F�l�D�?9���2�La��0l8A@�.`�����~D�+�A�7��L,���03%�W����PD*,� V�zl�4����do�$#(��U�����qp�Gt��)�a�n�黜t=S� ���5q}Նxi�mnQ��=���~�. �(H�=�H����S�[�v._�y�$�����Z�󜭗aZ��{���KeR�4^:�����J�d��3h�2~�PN��'�)v!
��aF$�(ᜠ��8�r�A䭸q��Ge1��&���5�c�d�\����@>�ӄ��O���tV� D��xWY�X�[(/[�bIA�%��������0�JK���)v~&|h��`:V��K��2O��g���MˈD��R����f���T�>w�$�4k��
�@I&��A/ #=�$Jy�S�s���o�s�Q��;�����y����%̿�)��h&� ,�> Ј�aW����{�O��Q��%�E�9��`��K7N���j!�yO���o�5��8VR ���KH�o,��b��+Ҽ��j=b^��ר��P��,!3�R= |�J�"/�{����'��>{P!����Ks��?�\1���(W��=Ux��Ҽ��0�6".Q��X��h�	@�v'�X����=��Ί���o���ePT�6��qb,�e�LQ��!:��`�Rzb��zz�.*��f'��{����z��)�a�m,CM�@���"��"�V��5(�O�Ā7�i~���`_Kc{ ����};K�k��}g M�S�҈����?�����M�R�ψ@e��W��9{A.�+�!֓k1k��a�J�:�&���!l`�X�Q�n
�&�w<�Z"r�VX�aԇ6HL�gׄ��2=N-H��$�'�Y�^[���F�7Ua}�f��Y.�܃A �a֡3�_�U@�1o"	O�(�s��$��47��'n���$��F��#�ex�CqL*.70��F�s�Γl&��y�ԛ�XX�[q��5E��|U�!g:�SE��JLR�	'us)*��!d�en_���.��q��K �������a������1q�~>��tso���! ����9oQ��p�"�X�:MP~M��A����xWL��YX�q�
�4P�'��Ӟ���7}��~}:bw��zZ���zW������|\��ށ��J��ۣC�V3;G/��^bd{BfT�����"�ga�����)[[�C9�DuO�*t5n�4q��vĄ��F2������%�:�uc��'&?���V�t�D��J	U�ekI�{�mR�"����+a>�����J���hR��v����u٤	ȔtZ�tJ1P�Z�ի�+¼#I/�~�
�	��0s�����LV�	Ŝ��J�J��}L��!��L��uU5 @��������Uy/^����@"�p��tK�[�r!a�@��jaTp�A�D�������Pdtb����n	�w�K����E�Ob���y"\-��iW��:�i�.L��N��zlS*��e�U��ZU�fP�<����ǃ`j�e��-����?'�����֘��r���R������Z�L��>X���k��<�=�]�R0)d��oo0z�"�h�y��{�R�I���}�I]%
j�1/�i���6q��:}\j�ߙ'o4�;�e,�,�V%����5�|��Fv�Mw�?k:N1�!g5��anڣ2�a�F^%�ű�����V�����3�
7���v�eF�X�k=�Ϡ$�Y�U*�˿!��0B��B�����q@�k,��7�0[�t�@�@_��Ĥ�ٖ�9Ϲ1���S��ZZ���%I��S�c�PI�{��_��q��w�.Q{$Ա���-PHĤ�R�4��":��~�wp샏(�7d~��y��S�~��燇��X��Nv��o+>��#�7�6|ԇ�C�Uq�	2?C�)�y�J���������]ϮѦ4�b 42�q?��>��;~����`|r=V�T�i���`��W� �o�� a�m�ma3)BJ�+�������Ĭ>�Ik]�k03kxX��%3%��DB�]":/��Z#L:���,���?#���'B����m
�#
x��1%t�Bԝ���vly�_�7�'V��>#����yv�W�L�c�E�U�oF�}����SԷ��"%CO�\���k���f� ����e�����8�!d!�<?'�b���)�s'�z�y1���a�Z��J�4�ܳ6�B\�t�ϊ�B�1x>�J�J�1�~�N�Z�5+ݘ��5е�X��j����bf&��e�TC5����+품h�gUne���r�������(F�"vz7�f+6�����۠�Z��l	�;2[��I����X��,ٔ.~e�wf��r���&DXF�q]�����K"s~L9r��z�����!�`�?�| T���6��&���pX{�����>�"�&��F��
��>��V�b�ҭB�|���=��]��!V�������%�P�S�I����O!����?�?���SA{�I�����Ö�������b#�BP����fS.lO�%SW��L�1�j�m�[����7F�%y��Q�^��SǍݗBp�����Ț@���%T���R�Ilf���ei��̊r`��%��{�7N��X-���4M���F�*.�vSJZCc�A����1��S�����GX�&���l���%�fV����!��U��Ű«�T����G�e'>A˖��"ٗ��:9 �(�}�_�ٜ�N�'X��c-|���� _ReL�&�&�7�,���'���1��C�ď%}� �:����g�X=e�����@�iR��z5=.J�a�R�6�Dq��)R^��e}y��N�K@�[�sĄ<	�+2 c�8`����+lwC���6�m�yQ�j� (h����<��TqbN*V��%���}aÇb�]/��\��Ux0J.'F��[�����x&������J_�U��&c�D�ݼ�s��?����:��>Q.���XN'@@ԣl�OA��3�"�.��m��@b6G�oxmomw���Y���s2���(� (`Ĥ�����Z�/g�D^|`��N��^��ʐ��zZ��e��ON�����u�f��mM7?r擪,!��8����,�YJ"��mb�V��1yy��A�1v��Y̩��laF�LA�9bG�b�E��Ӱ��j�Yĥ듁1)b���*���I�5�(��xk�b�L��>�R9�>�H� �\� �0�9�g&D8a�����+��\��,-wB�f�HȔ$ǋĞ��b�F/2�_AG��?�C��~ԡ�v��V�7\�lr:<��V4n,
�u�ǤP�&�o����̽���<���U��r7�<[7$V��0�_?��`�ط�nWV���d���Y����?Ji��dt_�W19SaR���.��u3�d�kWδr���'�� C@���|�\L�1�`����rQv�Ӳ3Pt�J��m�S���{4�� %o�.�VQ:��Ã�ix��<Ν��ʕ.0��گn���n�3̝�a:���F��s%"���(����OHD#1��K|4����?R A'0"a�	��s�h��)H��b	>���A0'$$& �Vt�F�ۺ������8t�N^<����ak�N�;����.�Љ�s�}�OP��a1v�����yd����6)-��Q-]r.�	������5Џ��������?��g )'ԼM��k`j@nCS#�701���.4F�^���h�t 1�&�ڴ!��������龴�^uU� �)*I��*�wt<���c�_�UKѡ�A��U�&j֮��uy��X�]�j����gԪ�Wԫ[JM��G���տ�H��7b���5,�M�s��g�SKC��0��N���
�&�cmJ���Jݿ�o#lȣm@9\�!:�s�5WX8�.8�!�J(������%^���S�?c���/ۋ�3�ah{�Y���z�(8	;�!8�	�Ǝń�0n�d��2�gLC�͸�{9�/!��<2rO�!��sw�s�,8��[�z���b�~��؇+׏�j�I��:�,:�|�!\�9H*� ���M�����Ϗ$~��.=��L�(
�܋2��$v�B���T�|��~Z��+V�������x��@p�+7l>��q	2��æM���\�5q��!d睢9=�����ذ�;� 2>����w	�o�ƥ죤p.|2PX~Y���K(�sw�\GV�iܼw���y��q�GV�flHv���NTp�Bw�^`b
-+�� �4S���U��u�����AhH��Ev�H���$Ry��u���	�o&�QT&ȄS92����P"�H�Y�������m���{7�<Lj'i�����49��݇v`�MعoҎ�ľ��p�J6�>~B_�]�\ޏ��y�4�Σ��r�L�Maj�3]jC�P�#}-��T0���kh� ���T8k�z:V���ym:CȌ�enc[KX�Y��Ί֙��܄�dH�ҡ�\C�Yu���Hu��c�q&�7+,jC�Ѐ@�O��KS]1�)���>@ቄ��ѵi%�+$�Sęr��dըU��j�^�g�P��_�կ�M�w��0��jaa+[3Xښ����̭�3���Ϣ����5o
V�-�����Ѷ7�ڊ=G�cǁT�߾����$'�1����C0"�'�T����°�����B�6?�������K��p��7=��0�t�ݐ1�0s>FO�+�A4b(F�K�m�M��	�~��t�ې�O
�PN�E\�y��t��4�u�e�I-]!��K9G��v��Ws�鹺H�:O��@��SPGϧ"�*}Y7/��n�x�^F�Y<0�盞{~�E9@3�}J�$^�˪i��Xuۿ��({El�d�sm�%�}|����y�Z*�W�m�R�v_�5^Kq��N��Ɖs;q��n���G���7"~[��S��K��	[���@m�"5��çדrHckq�D��Ş�aؖ����%1k#�p�rL�>�����K0y��.�Ƥ��0~�h��=�j��i�Q�=w:V�XJ��j�?a���^���"��'�Pm8A<�!vPX\"�ew)t�[�#i�l9����!��q��I:s�O��;�3m���Ŗ=�p0�����3gQPR��o��Ai&�&��c�N���~�#�8ɂj�f�06�:�$=�OP�=�t-��F��3 �ЌH%���1$�hL�1��@k88$56�����@[�N��̨F]{uCGn��əw�,�}�rr� RB�057���)sX�Y
7%8蒪c��!AN���>ѵnۺb�S�qߡz�V]������,�;A�A�v�А ԤQ�j�����TА�p�$F%�hKnC�`c-1~��@L�=	��ͅ�����D��BtR,��ݎ�G�cW�n1��si=b���!����M*��ڪRB�
(���F*� �p�@��� x�z� ��Ҟ�`)�-�1����@'9CƎ���<��'ǘ��1z�h��8S�M��m��}�2n�࿷ΈAQ3JN�2U�n<����q�`�]|�2O���t\�q���i���Z�?�Ki��yy7��R?@P�J��b=���n��}[��w��p�C:_:A��w�&9:R�+V���	"a�`�2���� z�����؉}R@�K��� z�����D�\�<�}���P�F?��8����ݺ���'q��a����փ۱i�Vlط[o��#۰��&l<��l@��x��G��8�
�i�؝�{��a�MX�!�j���� ��[��&b踁pe���2�#F�L*�fϛ� � 8����/R8�ݴ	��DM9,�����d:
�6��A
g�l?t�O�����8y���;F�>l�yc���JBJj2��݊��!��i�=r��]��w��u2/ѽ'�aղ	�<�����KR*�z06у!È�a�	H��WN���}x_*���X:����Rv������pI�ߘ9vF�I��08�{! �[[�y�IYi�Gߞ����"ݛۏ4Я?).RC�&Ftϖ�u�! 8Ñ�mcO0�$ K	�f$%?t��A�!:ΠcE�YsRx�~��g�T�'���ϨU�gԭ�5�����G�V�a@�n��2��1�7i$F�u��a�!�t}3/'�������9w
������@�oH@,�s���BjhAhs�V1�J�M�6#is2bVb�x��U'�"�I-��2� �3��E�Η��jȗ��K�F%�����Gp \Ə�!}g��a��S������:e�;a��a�L�٭��E�;�*/�
�/�f�%�*�����m�G��ɿ��9�.gp�''d��(8��9��q�$rn_ U~��O�b�a�ؽ���KG���ً�қT���8aA0��	��b�m�� ������_����Oj��g��  ��C�>� o�y#*.!��]��U�M �{`-�߆+��p����2�W����|�2���q�GXxV�R:��|\/���7O#=�.g��I�~|H8|D�P�'�n"��#Ǔ	H��X�z4&�
�1pf�A�T��� cL�6
N.��҂�	D1����Z�?��}���$mI�z��KI;�u�nl۽;����GH�B�ك8v��t4[woD�D�IS�F�ux��#H=|���q��<���|��P����qp_�B�a���;~0��\xRaneE��D�+#m���rڦo�ކCoB�227�AA( ���#]o(��F��8L�6��O�$�}��2�'�@beĪH���mL��x����1@����+,�,����`���p*@y`�a��*������Ҍ�_����:�Q���84�	��s��X�R�Ԩ�������hР7���5D[�F��H�7~���IS�`�*ȇ��u�0���);r�ńɣ1o�L��\���(ld�C����8�۴�����Fڱo'v�E�ظc��O �^'��"BEJv`8�(���&8 >A��P�xi����JC)��؞c�q��=�E���##S�&��t���{����8gL�3Q�o�,�@iY�n]Di�5�,ܾ����
�������v��#@�^��'�q��~�
ґ]��[�ϑzOº���r�v��b߁$dd����4į'@�R%���"q��^�{zO�cLʜ�����޽� �5|�]��=	��"��6��x����G`����#$*���*dAc`�?��|����Ԭ'&L�����ػ'���Ů�k�vt3�_�G��2����K���ݳxz���?�����vq#��؂K�Px�(?<��w�F�:�9�#���m�+"�c��DLY<�����
�V\��Z��f�	]t���/F�ncC���A� ���@�!Ga�v�ۮ- 	B�� ������/}ۃ�GRI����=��igj�eO
�g)��H=r��yR����U9^},BN�>��x��o>��9�CF��aBT���Z���@
�U��pT�t�1|�	>�3�4��n��vB1T��g줱�0u<�ϙ�Y�gb����0c�L�9YlLʆ� �ᾞ�z�N��59��@��l��
r&5r�p��6n�(�w��,��Y���2��h��pWo:�ֻ[�.hױ����H�ԩ/%(Ԩ��ZB!ի_H-�~E��I�hٴ� Q�^]0���''�3��`:i�����9]ӈ��C �s}RL�H���%���X�xlܙBΠ�����T������ز{3��Mذ��w�zD'Ɠ*��-)#�@�0)��('.��!����)�ԑ?<��r�q)�H�xk��a��	0�7&��zM,�ae=���4�G:��s��y� ��gQRz���e�(�_���P��`�*kw8w�7���f:JK������Sri��1s�\��"4x�l
�g2��'cӖx�H�&�z���_"'��b}/�.�Ɲ;�x�
�} %�j��G����G��n��KV?$��ɡ��x���o����=�M�"�
�����b�"K(�U������bނq���p��0�S�"8h>R6�Ɓ!8|8��#q�LΞO �ǹ�	�8{!�O�� �uw(v����86N���!o��Z��)�1kָ`�,��4�� ���h=��ӛ`�K���a�&��e[L�5		TS�BhB8�c��ꇠ(?x��7���"�ې�m6n�I�+���;��Dj�6�9��j����v`�ͤ�RV�h�vھ��a��Cز��S�n�������/������Ò��1q�3���#@�`�ȁ
"VDfz02֕Ԑ�j�Q���؇�+!�A�ۂ�H�0�]�>5�	�gL�L*��.���K�b���b�˳�3�&a��:�9H͘�u�,<=Rkf&���&4��s�H̚;�����a��I�2},&N!(�u��3�v�hAC���y��^�ڣZ�kA��!��]�&A��Ȝc�T�C�5�@�+M�5i����g����0Ę�C	B0w�T���HP�����H^�&�r�� '{RƓ�gb�j����M;R*<a}�nL�*�7��H�-رwM������6��ZK�*<�gTFrz����c�5!���t�h�q�ꇐ�@x���w	��c��Y�2w,�O��a���2���ah�$F�7�1���B�j�.<zr���C��={z�_�����:��Ww����8~('Ǣ(� ��lÑ��
����-1tp_�nJJ|8<�LGp�b��y#<���+��A�>K�
Z���D���)ȸvo߳��]�*W���_D ����>�K��އm��!\������]M�?���h���9���{�x.���u1��Y?����:6A�εaj��ic������Mː����D!�L���Eډ�=I�z8��Ec������nز~1�bfc�B[,�i�Y�1q�>\�j�ʢA���>}yT�hѪ%�Z�6��� E���k������i��Ts��# �1��Up�]o���oHD���X��a��`���m#(n��م���Rm2�vo�6.�R7�:�I��l߻�j�	H'p9���~�W���η+Vsɉj�Th�c�p[*$�aK��)3Sq���Kg��3��e�m!S�3�2�����`;����"�ܘ�c0u���.���+bɪEX�r!,��9gb��ɴ�H�H簠s�C�P:S�L#�9㸍��M"u5w�L�[4���.�.�ɴ��0v���8����)AL_��@*EC�7��ꌶ~G��Ѡq�C��!�W�H��� �+����֩5̌�1l��uf"��C�����a0}���j��wVe�ǎ"h��������R�I)	�B�h'g��uHa��q�#�۵o;v��EW����JC��O��h�~${̺8�.P��R8<���W�%�2o��Wa������í1f�0,q[�5��\C�0c�+�3�A0ģu�aβ���
��+됗����#�U�Gc�ZW�xN�Ϫ�������󘄅sb�$SL�h��3�|�x�X2+O��USI��o���JX��C��'����(���ȘH�%�Q%�^�zN����������c�o���+�!��A�H���m��Ra�+Wτ���Qz��!����'�!7�����6r��Ĭ?)�����M@��T�t���5E����P�;�,`�P�v6��a��8�SFY`�c�s�ǈ�Zp��K����C��w�.M��BϤzkv����t턶�[S-�	~�U?�n���c��X�	{�Aj.� ꃐ(�F{!,ʓ
7�p_�y�戚l��-ذ}6�܎��Խ[�g�&�=���vb���ش�j��7Qa�]�)��ڲk�Ϟ��{��>GI��O����R�$F��i���;9�b�`�)K����* dB�!7" ��C��C�n����)VD<�͸�cE�mƜ�B1�X,s]L�h)�i�4c�LEJ�	6�`L��g�]#R�氵����A"7��7u�D:�d̚7sLÜ�S%�'�F�q��A��6V(���tF��x�on/j����<�i}�P]�Q��P���HY%q��ߛ���-��3L�`6�ќ����I>��9N.����es���p[�}o�p�(T��ų��m	|��N���xlO�T�;�l���V�&��
xO�n��M0�|�]l� ���'�B�' �H#Nh�g#������un>��`�,L�=
�a�X�9c���X{RDN��t*7z����:�C#������x����5����6x���=s>�� 1��Z�mߊ�Tyڱ�*RQ���"��^ �%��\� ��&�q����Eq������j?Wx�ѳ��8��%�$#������f�-�|����܅�s�`�Xuۿ�B����˗p��~�J����(���`�^*l��t�T,��:�jOAa#R^T�t�ZE�*,]9�
��H5=.h5uy8����tu��@�j�4{@���舾�:�oߎ�׷�kt�&{��г4�t��������r����֕�{�w@�n��Q�k���G-*��4�B�Sw��7��� ��8����M����Gy ,ҕ>�
�y-���j��whs�l!ߚ���&��ؕD
h36�6nوT��l�H@ڂ�[	\۶��ۍK��P� ��\ǹ���j�N>�
��V�B B�H�����)�GdV5�*� n"��8�/�Ch�p'���}h��q�6{�PD������B��V��p�:{&LK�h�x��� K�X�{�H��wnjnL�Ɯ
{��0v�(�;�%�3�����B0�JP����c�d)��e�#�`Kp��]RX�߯:um�Vm��i��R��>'.HC�pQ}���z�hݢ	����4G���`i�K��c'9a��at��� k{N)7%%dFߕU\���>r�H�f-��Ϳو�`lؔ�-��c+���7	q�u����{(�:�gw��݂M�6����-�D����fܟȟԏ�H�
�:"IJ�a�8�3�O���.p�J��PSf�I�F
��&t*���!i�/v_�CW��\�k_AF�\*8���'p���9�i�w#3�,J���ٛ�x���n�VI�]:B�e-����\�@zV�	B��K�|:)%'t0���!�=��3��@w�����o�P�2ė>S(R��<���`����D�c�����#�d�S@����@�w���ɣػw/�Qa�k7��R|���6o����B�~��a�τ��b�!'Y���<���Tv��9grQM�X}59��t�ٗ�M}��-Ch����&���ӡ���fF��h�7:�ҧ���>M�EN�0٫w7���];�NSc����4��~k��͛�֭�����qfו6z�f��݌`&A�$@� "DΑ�9��9�s�s�V'eY�J�lْ�d{fd{���<{<�e�u�:�bS-�j��y�i_V?��J,T}a�{��>N^��GbF&��z������E\��m��hz*�S�}�P���������z��C���u<~|��­wMϲ��n���wq��*�����7Td�)��w~���/�7��&>D_�%��$�'#�0�QJ�%}$5����C�@�� |� ��H�t��q�Ó�d*�Rߥ���r:�J���^�ur�I'�C)5�FET����Trq��E�H]Bx,C���2���<��� *GS�Q����*���*�ԗ����%��9=��mDt�����^tNpt�����D�����M����mh{M՜%5�'�x�O�a��ꈰpo����T4����+�D:!�t`r*�ɉ�������RJC9_C�ƕMI���[�u�A��(��o�5��mڛ�z����c�y^�x�A��̘��&��:���9*�ySĳ�u��z�:��/?w��\d�����D&�#$��=;�`JF�X�6+���7�ŝ����g��l�_��/}�.�-|�w��gn⣟���|i��ͻ�O���,��+_��_��&>����^���&mEi��V45"?7�!^��wC|B�4,�Lbau3K3��4���3T]�������T����dZ`�� ���O�^�����o@����g�>��O����TCo1ʿ����_.���}d���U�((�Gee6:y"�љ����� P-#�RF�)��'T����s���q�,�|��UH �Əe�mI1��9Qq���Ep�7i~!�����^��|/��/�B�����g�|�N9�	[�;�ĩ3�pp=�Sn���Dtr:j[:1����p�[����������ct���Q8�nޞ�ZZĵ��p��5\���wVq��2n�\��[����p��n>��[�kw4�h��>~���+#�>���
��~f��8Y1��',萒h�GR*'�#)����:��"�  �x(�J/QQ�)ӖzD�̼L�^�1%�QS��r�f��� �c�  	Dm�M�m�DqEr.e )#1��6��$��L������2�:Щn}���o"���S
���B���"��,]�pD2��1������ �ت���U ڷol����C68|p��G�1"��ps>���n>�ΏG��L~�|�U��,�6�OL�NIFtL,�#�L9yna��JL
���#����6籩95��p��U<|���~O޺�����]<z��q^��;O�a����0�Le�5C1���%�nnF�fN����|=`�x��<�	�����=��pwx���O�	�gb`�W����1<|<�`p	���>��e�po~zo���������G?=��?9G�>�Wߚa�4M������.6���OBn�?B�>>g"DE��"���1�ɥ9�h�4Ah|v��q�>y�A�ֺ�&�_��g���{����0z��5��-�t2X�g�~����;���>��>�*�|�-����p�>#:*�ҒH���`��mlޞ2q�����2N3==e�����10ԅ�^3^P���sR��r��"ʨ���p����e$��f&J�S�̠|�2�#4�!��	"p����<����zRyJ|���Ϝ�I:�㎶�s��i�3p�v�7����TT�ՠx��m33��FI!��E�q=��?�=^�nFޞ�>�f������̯Mbys��ַxj��t����I��E�nЉi���U:�W�_�C�6��Q���ԴP:�(�B ��Ŵ8�J��L$L.*-GF�D�K�.��(^�q��	i������DB(i٩O-�0�T/�E��-7Us�*X�����@�����Qy��������@��0*�h����栬��(��.��]�-F��h�$�Zk�Tҝ[�a�m4�52Fsթ��T�TD���p䘖����s����Cۍ���� �t���;z'm����[\r��ĥ�T�Ҋ���R-����<�T�1�����Z:��7ԁɹa�-O�T��2��^�M*�{��0���v�}�5>�m�XB�`�G;01;���)�l�P9,�6QWo�$T�3x�����q�8�C���v�糗9�}]q!���g	Jwd�D��!��04r��Ӂ����G�7Gq�� ���z4@�2���{=<�p�V�n�bh����W�s�' #��՗�+����0 @um��>�Ncjvs������u�̏cmcw���9���O�`imW�p�����7�����{b�Z�����������h��B����̧������J���l��"A��90wb��z�V�б&��Cp��i���j�RS_��F�e*��	�i�I�M�F8UO��v����w~!~8��h�<���RϞR9Ƽp��g���P��z�srw������q���3��?�sn���?2�p�r>�+��Z���T�e#3%�~.p������N����������������6�����(��AF�c��
�\����~sW�/�"�������{��ʵ�/����
��3͠y��X������R����1 �|,
Q��jz��3�A�s_&С����F`$(�q��IAF��rQN
�AT�kJ�+�tj����Vg�I4����D�4����ۻ��RY)�����˿M�A�Md�̡�+�d
�k��k��2U�U�	V���I�w��T���@�!<J� M�T�J��N���a��7�ٻ����{�����}�`{� ��ɣG������������ru!�J.�哒!XS�Dq�G��H'��xnTի��
������&4Y{q��@�� ���S p�����_ã��`fa�|v]C�7]\���"Į�ac�*�7��:Ͽ6���8fw�	\~oA�����a��a�����~�.G�`	��f,oub�z֮wPy5�q#6�5a�JV��	�F��Z�V��d��%"#S�M ��|������eЪ���ު"�$��؆F��aLLO�\�!�h����9=����4j	y���Ƶ�wx��60ڠ���o}����N�����Y3pz�����ۿiE������o�co��W_O�"�^}�;����eF��\����p��½Wq����k�Ps	YI�!ʡ(���c�㸋Q�J��X��-N(��15;�D횟KG}1�X\2?+�N6�7��WQx�??ۏ��q%5���<ǿw>Ї�#J_�]@db8�2b��s�%�t�����HB���gO����th/a���;>��]/��=�h{����7�Z�0:3���1LB�tLSKS�U� :���X]����(�y��O�0z�@o����J\��Czf,��z��^q�vS:�
 �=V�K�>*B��)^l*x�1I'|� �"}Dt�5����oQ1A�)*�(B���@H�>
�֊��S���,�b�b����oKCAQ��G���ʚ2B�Uuڪz�R� ��<((�Av~�鸠�b�7�N����'4����
� :��ڿ�����8q� :v'	0�'�Y��1Ȼ��l3�H�Ӳ4�HEߊ&��y&��,��ss%�:��AU8H5?<ч1ij~��H+<�k�U�[k���*���G0K�x�� 8��EYt�XX� ����̂|�[����/c̤d/M+8�%0���1�p�3+�
F�<�cR��	��b�t1��
�Xš�*��(�V��8���!�
0�qo�[0ϣ�	��7��=oh^�|�8F�LzU���mJݩhc� ��p?�e�ga�'���h7���155��(_��e����T��y�
!��ŵy�_[�/���Y� �W����~�����|�<|� ����{�_��׮��#F�s�t�8ʋ|�ѓM)��7q����X+�j�W�A'�*(�S	�̗c�i6�T���R!��*���(U���Trz���4:c��X���EM8#�PB�0�D!,���4�/��P?Sy�����h:�� FJay(Np:��o���?~��Dm��Ǒ{��v�f�|pǇ�����Νxy�^B0�]���1N��w����\�b�vF��0�����MU�J�^�X�(3��&�邋"͙�>�raO�cM��L��Q*�mA/�d�ilH=�T5�ɬJ�]"����"U�5�Q����8� ����d:+�R�|"�X(&.� I�R�S���m���HEb��ʫ���	F
H,��iA�/QSk.�i�V�z��	D���DTC�=At��Ȗ����c��v�������H6%��R�B�Ҡ��g��)1T�ɸT�gQQc[-�;���߆��J���*�aLR�H3+�T!�:�<���~�X^����	9jO/g$����.6���������UͿ��c�1R�N8����8�p�@����g9଻�Y�R%������Ho��"�}s�<�8_�&�GT���@X�B"��L��:l�p֍���w�^s�����9�o�DM2�1��S�v���R&g�\��~/��kQ�s���weeA^TRި�/Ń'wp��U*2M�b�K,o���~�w�������3������+<�0B��?����'?�����?�'���ѽ�6p�v7�C��z;���WT&��&y��;��0׃��B�JE`щ-G)��$���R0zM�SN �N@NA-X� 2�2���sIt 	��F�iy�&�<��ƅ�j)�<�H�&Zsm�X��X*��}����y)Gp�n?��>v�̪���0�bh�
���;��+/Dƿ���W^��9����
�-���@KO��;�7:���a�O����.��@-fj��+4(�J�
6�'�Z$H�� <�RL� d d��4���ҢJ��"AHcC�PQyJ!MR�j�0���S���[�&��r��2����nꨭ�g���x)�m%���d�䩻B>ac��QM�e�M��
�7U�UVY�b~�TQ&����@�������%�*:~²P��q���S���q�10:LUt� 
���A9��:�>cO'֜�3�sL����*(>Q�C�TR����Q��f�a[=����݌��Vt�k���8�3���������GM'�������j�"I�8�� ݃'��!��O��`zAU�TK��l!��yM�=������Ngp���'b>�r�f\7ϳ8w�~��s�4VJ��aԓ.?W���9��
�����$���Y�ɕ��}އ�P�	ã͵VX�m��R5��������S�c@�y���DCC�������r�9����^�{rkWW��ݍ�71�����5��׿��'�{|����r�7	�?����O}����'x���D7_�#����hC��r����x\j�C����}�7�16ڀ�Vˤ�T*"�HN%Tm���|.x�yCU\�g���#2�V� �t�S
�JG�&0��O�X��	�� � ^x���$�)&.̼����&йD��{�*��������a��c;v쐙�bCg�{�n�ڽ���{�bϾ}�KTC;p� %3Y����Q�LG�Մ2^��T��7v��w�˔�к�[�*jPU'%�oJ�����2�3 ���o�z#��%یє��޷��;%�ԧ@�M�ZP���39UcC�t&r�M��h���Q��`$u�1-"w��I�(U-�R�����gQA�QD��Rscj��hn�EK{Z;��Q����(E�����}�{�狻��QEсg@dY�"�"��tm��l��)�V��Q���̼��`��g<W�*;�*[s�.�Ě}�KH��R��@���+i�����h�&����*�R�����,�ߤ�#��a��+�ٷ�좺9Ġ�I��6��j��Wo�ۋ��x��x}�ө����98�����+��i�vr�����>�r20q1ci27Og��ST�pvw��YG�>{�n�p����R_EwoOx����y���[�
��y�D3H�q�6���͕f���Ǭ��� J�u�	{�N�5>>�c�X]����i���AZn,V�������r�*�����g�qe�񛿁��P��g/n���oD������������o����Ǐ��G��(om���c�xr�9_@��N��L�of�蓼�1���F������g��Ѕn`D$���_���j�	L���]��?��@���C�p�4Y������X]}p�ܝN��K���8��n�����r�n�8�r��=�l����8y�vǎ��*��@�Nˆ�Ѭ�]��2a���_¿7J�%��CRzR3N��䠴�2��榘"����4љ��ҩ��	�t�������@��5Y�t����]����1�H ��Rϸkӣ"��)śԜ� (=�1��L�,U�Oǅ�l��G�Ashں4��Yo�`��<St���J�'��Q�DZ�!:6��C��
 R�W�k:,XՐ�,4�՚rn��i��jj�3��V���ҳ�M �1�s���N�L�jw�րhA�wD2{v�|j6<~��m��WP��^��ὰ?ùMA��I�3�;���3�+�/K�����*j�Ԯ�ǷgpD۪��J�k�����8:���g)�x�����N�w����{8�����t�>t�	(�*@m�e�]�6]*v��t���,�����	3Km���Z
�}?BK�v%��P�NTKn�^Ƽ���Os��CH�т��nd(��o4ϭ�:Wb�bW���2§�L�Ȼ�n���q;�������|���B������(��k	Ȱ�h���7b��m̯ob��-\�u�+��v���}�����|������D��37=��|_�կ�������>��מ�p���~����br�Q���q7Dgסg�F�&1���_��/�3����J�d��	�
I���O!aI��	DJ�����R�{�;c���q����Icx�w%P\���}|����7��¨���qF�v2��YW��9;�ם]N��O9��SG�p��O��-��C�m�=���v�2�4m�#�v�û^��t`�Vs��#�= >���@f~!
ʊ�Y����D�0�.�\���Vt��=mt�u�[���e�ѹ%�ƣ�V}!؏Q�yx@^�=xAk��!��C�G�Y;j[�Z�i��T�2I �W����s��(�NVi9���^m}:َ�V�@��Ge�J+v�6e$E$U���t3�e���C#��B�EU�|Y9�|_�)����tTʭ�su�f��^|����iE�`�v?Rʊ�!���N���`s�
C*V�Y�a��m��M۳�0����v�z	����h��=8tt��]���l�C�����.�|MH�3�3�2LG�b�k�	�j��ј���u�Xk_u��`�A�h/���Z{Z�~*�:�TATm����
�燰��C�s����+8y� �z��9_^��1�L����T�SՉڷ�n�`.D熪'5g읊J�ͳ����x��=�1���j�"h����ޠH�O�Lr�c�<���4c���&u���)���=q ���38h���}� ���#rS[��ps��るTOW�]�����_�����zMZcs�~�!��o������:F/n�����30��~�?����7?�Q�{�w�{����TB7�Ǎ'�rw]M�8�Bs!��Ә��Y��¤Y�������P\�*>̴}�� k�\��	�U�+5��hUF��;.�	�Sp:C����us�~�`�}���yG�8��kUR��-�N;�0�ލNF���B��z����'�lO����ط����z'!�g7�V�]���c#���L�2|y���Ѩ�o bSQPZ���"��Q��Ϊ��m�h꠵7����N��R��C�i:��/� 
���^��LjN%����&u$�L3�m=BV����@�:���P{K圊
�>46$ R@��)')���6�C���n��jS�V��J���K��j�rȔqGIe�f!� �J˕���*.AH)K�9tx�T_m�Mtb�?"U����":�cxʴ�9�}G`/A�� �Ɖ�l�{/��l�.��I��C8�#���{��lL��S�U}���<� �[�q���W�@TDE�f�U<����hhm�w%�;5���AG;A�N�������Q��7���jB�����/��/��I���A����{߇p��.��O������5��M@Q������'H�-2�uuY�Kz;42��\0�=,zB�xBy�JZ1D��Uz�ZH�&���M ��s�u2���I��ۃö6��;�y9��V��S3������
��'f�o�q��l��}Y�R���a�����*�k��"��+��?��������kQ���r{��hF������e�{j�(}�1�>����w��`[wP^�
/�`�Mc`qӨ��������w14T����\���"gh�.>RB稂����Q]v�Q�Ѷ��?�ȗpq��1��(�ur9���!��X��)o=|�1ݷ?E�}ZT��b��w���'����c8v�(�ُ�;�۷�@"�^ޡ��nF�q�����B�a{���Փ����G~I�

PX^�ʆ*4<�[���A%$��qi��Rd� �tn����V"?:_�J�G��}�YՑ@d���
�Ht(�8����gSu��a��k�$E�1���"T7T�;עUJ�jH�SzQK7ԙqu�.��RA�Rg1�$�4�(4��V1�Ƌ"�H] ��okΘ���n�w��b�;]Zb���(#�Ț���������ѱ��!���q#�"��l�}ۓ\��1�Z:Bk�s�u�����9u��Igi�k_KUhb�V�M�N�2�3�U����yL�P`}�`�L�����2*�ZL�����6�*6�t��=���?�?�Ї/�L �~��{%��sn�+8xԆ0:bz�u?Oқ�?���R@aR�<~�$��/�*��L�N��5_ӕ��<�4)U��I��� A���(U�vJ.n��a�p���a^�GpB�G[^['������n���_�g'�2���h��ѩI�.����'θPy#.-+ׯb��L���S�����eL.�F�����&��=^��nOz5e�/n���oD�W����&�D�xw�x�_}��O���Ga��,F�*A)��X�v3��h�+@/Ʒ>��.��0�L@6���#�x���$)��r0'OS�8� dN��$�N;<�pvu1v��1=w��y������=j���Y� /�Z��z�)'G�ޣv�ב#8z� �ߏ�{��v�c�����9;N�I��;q���8��㤓��QѤ�]B^Q)r��PV]��NF�C��֏��>���3��ct\^B`D�i�Mb�O'}�
�|�?|"o��/����e��Ve�����t25�UE�5]g��%��n��F�?6nDg�	Â�:,X@���J-��B�
S)'����>k���/���2�#HX��D!6^i�H�Df-��X�(���ʚoƈ���D}���,���ʢ��.h��v��RΞޮF!���9�@� !���H6Z�UՎ�U�H;��Jי�?���?dcL��
"�3�Nf�����z\���1�ȡ**d`�yO����4ʨ���*��-�gmTCm�m�CQER�S���`��CM]%��N��_���K)�W>�W�����N�$)&�5Mb��?��u�ߋj�Ł���b�TͦJ��A2��1���
a���9sm�)��F�vORJ�U�B�T���D���!,]�ꦞ~'	����up�d&N�q'u(�U�'���"� ˴�R�(������,�f�����'��a��&&V1����+�эM��&�f����՟=UC/@��o�&@���_��_ƽG��F�"|�>���=��^��ǫ��/�OH �
+0:����y�,���(�Z��g��+7���y���� �5Z�}9F������}M����g=���T��M'�Gՠ�?�澞sru����iZ����z�eG�r�ݝ��␳�}_��;w������Ýps>�THG��0���C;���l�� �ھ��p��;y
g��]*��3jBYU*�Z��:�3�O���z��Ձ�:��e���Alr"�蠃�"j��0����%�Ǻ*�"h=�2����#+������YӾ��Lf�3
�10�2�Ht�
�V�	Dj�c��N�fi5�5T��-�3��W��m�(!1�t|PJN�9�EFN��dde�Ԝ���ҏ���,����.�ˤ� Rq��ۆ�9U�!Z��N����CvGqHʘ���1$Ja�A iy#u���1=`���(h;'�9�Κ��/7�ȇ�#����##Y�j��\1ʫ/�FYA��AE�9e�-h�n��
d���7�Ǆ#(,� �B6�loo�;_"�>����^��!c;v���6J*m�Gm������3�+��]�T��yC�σ���֒��'�|��^����~V����ͩ�>�=(��<�.he]�o��"�QQ�Rߚä�;�)#ẽ�|<Mi���*&ӲґJ�gPVĠ���
C��aT7����??��ZX�����ULn,czs	�76�rs�W���:��+_6��� ��eͳ��}�71F�w�wf��zB�@����-F([���T�ڝE����\x*:�0���W�17׋��:�R<z��x��;܎���&���X�R,�t(�*9�@��yAi�&�&2ZO�Hg���^�U�@�_.GzN6���<����Y؞:�(�р�BH0�l2��f�45�����$�j$A��Fq��������UŴ6Z�SXA>�62TN����wo^�1�ۗ����6��F������������>�sQkw'�ۚ	�Z��b���"*!���G\J"�S�hE�GG#�h����t3.����($�����m��*��R�e�L�QTMr`��5�XEY��j���2��
k2�t\M�� ���B��9f�&3'�`��ͨZ��I�a��Ƈ��ȵ����_ʥ��+Ԛj9K�B�vj��(%� ҄Yk�Z���=GTzΑ���3��		R��8F�}̎�����a�Ȫ��||��!3I�:n'5I�b��4�<>8�dB,�ғ�~��3 )�~*��X�@�
5D'Rj��H7�7�oʩ��K
������G������Kp�b߱����>�����v���^*7�{��<�sP�q��=�t��(o��w�����J�
����;̓�;|5ǈם�>
r�O�ߓ�U����檅)���3Nq_8:��	H���Wy��{��-�Av@�x���MHNFVn�cr�300ٍ�!�!.5N��H)������61����eLm.S!�c��US�p��=��?�=�����/�H!����o�J�GНW��Ǹ�����#\�]{�U��X@M}��b�98�����[���T'Z�#�01���1�8���|�:G�H����<���j%��:8�2'��S��;�攎�b���T�2���*C/���J���#5%Q��C����r�l�s�p�8ٹHMO�"�4i.9wG� ;{F�tPJũi�����}tp�V�T�wp���'UF,kz�K�P�Є��^t��bhjC���@?/�ޡi�N�@��*jCa�"���KȾ�GR`,�� Y�J٥FqD8BT��M�w�2� \��	��ekS�[c!�Tn1Sn�`z�y�O@0�b�7��ԤTc"j����n&�V1�Wk���Ւ�K�&��f##[��%�Y�?h�J]�H}��T�R�Ji�՜|}v��Y�Xi��U��~s�S$���:�-�_cг�,*VPj��ő0"��L�a�:}ʀ��ñ�JkY�(�դ�P�Ä�1�kv'����;�83�!��dU�����l�0y"H�R�䢄 �j�G�
R��Z{��5ԏ�������5��(�
J!�}�o����#�������Ɔ ځ��{P�<��*pM���&�l�#�`{�8��H�x��3���9�f�TJ�pQښ�p��м"g�38�&��}��=�o�4g��w��z�3����Կ������i*"miT����/;w�A���.�"�*>(8�[�����l�ZXE#Sc���߆������W0����+[X�y˴��ML-/bqc���/��~����r{߂H�X�?}���K_�P���ȫ���!�BW=�"z�M��*Vn,1��1�exbK��M��������?,���_����ƭ5:�v3!*V�:�F)�SzEyhGB�AN���*��p��yѝ���鬪&: Ow'x�Y�,av��8O�iG��?r� l��������p"t��wN����s'ma���lq��a�߿��cT=��ÁCJ���w��)g:(^���8��H?9�]>��jQ�Չ��aLMaxz�3j�?�1n�&&�G@��g��J���H@jEUc-J*ː�H9����s�e!)#Q�1���7��>TmFt >�T�>8��k1Bɟ��B������p�X��s̝��2Wɚ��4�d�8�T���II����hk���*%|�^K�^���F�)�"H�Q}] H�BK:h\C]2T�)Z{HK0辺(X�)�+�&-Ŭ� F�����YB��u�XAt�PQ@c���9fK;n��@5E���vS3\:Z:���"���M��]T���U����жU57��t�����T�Q�� �G����]�ݎ��RAES�z�����wո�����/l������5V�������X&AI��@=�k�ށ��ў�]S��{zp�hʃ�<�qڙ*�����ũm 9(	@>�ޫ'��sNq_p���u=:��$Y�Y�#77�s�#w�'��y�+� ��A�oiiIf���L�h������Z�F@x8��c0����+��U ��r�Ji��k�__ŭ������w��������D���?�1�y� ��B�㪚>����?z��[��i.2%�S�+X��^�Z��x72���H�78
o|�sx����A������v"	#���HJ1(� ��NE�	]<t.�TJ�T�m�#'�����gq�[����0��oB��ξ�{pD�jy��:}.�sSaiEV�I:~�M�B��	�����Rt���	��Sή���頼͜���\��B^E9j:��l��?5��9ha����%���'�f��'12=F0�`��7:h�T�ֈ��˸ċ���4�pr����S� yXT�Q?��;G&��}��<��o�|��|�严 ��\-�O>z�'4�{A�"��U��ֱ(F����`��a�Gc{ W�u{r�?�f��x�m��ʬ�(��SUZ���*�U��҇OK���	�RBJǩ��ZY)%-�"���5�J��i��8����
W:p�G�yA<w�2MLO�J��q��(3*��BEcj[��64v���*�c��P�� �� z'��:�x�	%Y-a�M%��3tڇU,s��|��*�����<��ӄ�+A�N*`�<���}�����Mc5��7ڷ~<n���Y�P&�@��*����}����T�98�-e�L�jߝ8�-?Þj������ב�;X���#�U�J�"P���QY}٤c5�����3��fP6Du����83�u���h#��_]���:f7��6������y���~��~���D�W��~��f덇�p�����{X��=�ƽ�� �QV]���e�,/a�ڦ��&�b��G[� ����czi��M�_��Z��8A��*Ӡ��9s!)rs2�:G-`GC�8ё(�nJ5���#{*��5���>z�@k�Ziu+�Ҡ�/BE͖ԟ�I���Z@$i,����8/�ӌ�	!�s����؋HHg�^R�2Fy�}t6�b�7:?�ٵU̮�`��l����ms��OZ&b�p� ���=؋֞v�G��uKPw��RH��S��L�p���h��� :� S�-5d�7�b)l�rrW��դ�<1�>߼,��gM`z�y�|5��R�'�}�&���M��x��� Z�����f�P��L��*:�Lb&����|��~7K�b��j6g J�m��mм��te���ik\Cѿ��1wW7:�st�AT^����2cui��
p��%U�QD+��@A$�� ��
���ä�:y.��|�6���)�,�`��{�68;�f����LS�" �ҙ�?v���I_΂-��}t�~���$1	QT�)T���.i�ɭ�S��c��NUm�0����Z����.��Ϙ�_^o�
dx��ߩ�ᴳƞ��,ׇ�%�iK`4m��fO�	肘`�4���sf����Z��w!� ���q0J�O���A���8J�������-,_����ML>J�M*MG54���e�����/~���?� ��q{_�H���?��x��3 �v���S�?�+�n�o����H,b����QZ�gVJ��'l��K_�*>��/bx��,������]���i��3�W��H��.(����p�c�����s7#X���N���#D���M����"�s>�,9q: �Ni�ngo���y��B#��skg�c����4W�;@��/"13酗PR_���t2������8#�y^<s���<K[dt����ׯ`��:7�5����IBi|n�����7cH-��h�hF]K�����V2/+6pR	����FhT�I�I!�q��NOo/�[-)*
��I�@�
�.)*�g e}����ܻMNP��}}�e��i�xM��VS:�LX��jz^���}�mg�\"ݗ�t���Z�i>�:�[T�T�T ��7�[:o���� 
�ꌈ�5i8��
���('t.�V3H�Ey].�xT55�^�q�P� �g)!B�gtC�eP2�sbtq<��+���h�G��s|�]<`OuaK�q�0�@�w��t��&\.*''��B������de����d��8���TB��������W��n7'�Ҧ�w��P����ʯUe�I�R�R̂���YS�2u�B��^<���t�<n�9�t��(U^6�C�����a#����|����٫W1}�
����)pS���ZR������ � �{���A��o��7���#�$��޻m�U�G�9���Ә�]�,L�"m���� fV�0�4���F<��*�����_��?�����2�����UB)�ӌ|���CU����Vd���#X���c9W�E�E�J������q�����	�(�b���\�tya�|8?�Ii��f���	޷���x�8#T{�O��;Kg����$g�!����h��4��>BD����$��~�,mne��Y�Ҧ@���[װy�
�oX��Q`Zڠz��R�<5f�v�#��X��Z��@����LipCK��SAq!�s2�ZR�.0D�^��-����Q-1�>�C��-8���y�;/���zy8�6HAY�#��I	4�Z�cQ,��d��)(0E��F�S@�9�7��]�E��6hl,�~�����Y~�I��
`ٻP���U#O��y�\�b�.��s�<��@P�H��Z1M�/��z���ԡy@�c`�ފ��Է��Ai8�~)�a�ghj#3S�X����<��g0����΍�%�]����lEAy���T��'����ӓ�lU@�@���T#j�{��0�C<G���=�����4Y���*��.�2ו�\X'��A�ҳR�Jyj�^SK&��f��^!�P��_��o�hU�.�L�8��%�sb��}��^��T�m�?}T���� �7���K�&'�g109��6�J�����7n`�~c�j���!4� N����Y&b����G/@�s��� �ۿ�[|�_«o|7�����غsw�`����QEp��Gظw�������/�iL�Π{����������_������w�)F�-O/-�Ao5��ঀ$GzΏ��T���t >���3���;�|C�ǈL��0�=A�s����V�����tݷ��	�n����+/�3�Ш����d?P^ދТ����J@z~Jj�Q�ڎ��ntk�gB#�|���-bzeрHQ���*V�6�zu�7�b��U[B����J�c͗X\Wj��kv�0Fa�?<�^:�~�����0zx��9A��Y���:/��\$2�גQQ�GHX(Uf.�o�e�jx��Ry?�p�<���P2���*��� z�~���Q8��Bu�(]f}��&�XLc�.�U��@J7�2���I?6.����R����R��z@^�o��PA��gLb<���P�h���͝���M�;@���{h }=h�Z��S�H�ҡJ���NQ�2r_Ƭ��~F4���0A[�3):�+�6�x\5��}��Lh�1MH��l)u��J�1%�
�T�������;�׏
�<o�OO���U?S�+�]�����>=���i2�R����׿����1�&Ѫ����a�#�;e� M�y}Q)9KqR�E�F���ֹY]_���8�8��`�5�$�&Ƹ��Q��v]]���)����U��s+�FM--�1�%^K������������g��� �˿�K|�>�7�~ˀh��lFk��۷�L[10��-������r����*`�r1���!����!�r��y!�����~�]��?���0]��{LWa����e�K-�#%-�q1���"�B�G|Z�SK��@*#ٴ�l$f�!R�r����B�ʈ3���u~"M��>S���yF�r �Щm9�����P�ijn��F4v��ch=�&�?4oP�+�3�F'$5�}��N5D�hN0Z#�֩�6nl�\!�"m7nP)]۠zRJ�ꈟ-u4&�>��$��$���L�b�������m�$ �U��Rqr�r����ɦ�Ax����#<Rc�
ԵYcrRKJYz�*z�'*k�΢�踶�d�D�ϻ�(�9f&Inۏ=/e��ڻL�Z��+�����(�L�jl� :�g�_���DRu'e� � �t��n����qdj��}�sfLb|n�<70F���GZ��Ʀ���ht�e�<�JI/n�a��]�) ��� ��Ji�h��P��M�o���8F*�Vс*ߔNT���b�.��v����:N.'y�Je
���GBG�=� ��-������Y�SN*ZPš��;�v����������"Ӽ,;���M՞ҠR�R��1�k�G�p?	XuT���1q�i�Иp4S�OQ)����s��NNb��U�ImZ�s�׮a���	#U�	D:.�k+��/����{q{/��-�~����O�_���O}M^�s�n`��,ݼ��[4*��{��z�������M��3�WT��y~��|+�2���Z�h]�n�����/����;o�P7��
q���+���e0Z���Frz*�R.�bMDrV*��#�iN~i�)��'�2R��`��4�;����Q��L3#>��k|%%3S	�HPQ������B� ��~ށ��b�w.Q�5��_UPt$s�p�h���<�7��6�1����dac�2���)��ץ~��{
�� ɶn]���-Kb�~�Q��4&�i:�i:��¬���Ƨ'0Lu&0�1�f���ȴ���e���5K/h9!1�D�!tz�JM�Q���_�����Rd`Ru��T���mV�d?D?Ŕ�y�i����ˤ~,�����U��1�[(���m*vќ*�_R�=[u�NP�yV��U����xa���#t9:Eݳˋ&�����,F�L`��q�k�EA��ֺ���5+���+f+-0��*�{'��e��� ��h��P���l�幛���P!T�R�ϤJ�ؖ�ҔR�R;J]�R�=e��iI�Z�������'	MU�����@�h�Ț��Vﷴ�Q�`;�^)1�b<�iΎ8ɭ��ҟ���`�PS�9�ۚ�2
�5$��c�m�[�15~֧JB����۔h�Πg�p����"�#����
;��m)0X����O�����Ջ�Ϻ�oA��~�����_�*>�K�7�ܡ�$�ױH[Ж0Z�s����Pm=����QN)-�F5��U��0�:k���h�����A[W#���/ᣟx�,-<>5B����	�T���HJMA�*��4���i���D���sҐU���&�R�qbz���}1��'�2��_�3��ؤ8�Zx,�A�A���|M����b~��_ �C\j*.UV����c���آ�B�\cĻN�IǵEh\Y��UK;��-��F�*N�i�X��fƇ$-�|��u\�{��ݢ
�e�_�mݸ���U�9F�3��ܧt���,������4���FǇ���Įo�!�JPX���Y��u��������v���d��z#�L�N�/��' ��3��i*�Y�.$P��]�� H�g��Ic

dTf4/:g��U��Ԡ��<	1�eВ��n	R�.���ʧ���t�a�
shjԔ�@T>rt�tx3�����̔y�^��s�8�7�a��uK���>^S!
A�,IVRES�Iw��Ѵү&c��q]����`Yu%r�y�f 82>�<yn^��;':�ST�ܟ�\`O5#;��`��"���j���	����l�Rl������)Ok��>ˌ	��'̘�i�Ǖ
H)N�;���x*��F�n�1��B�����ǁ��a�h�� �1ԏ��6n����^!�f	�tNL�c|��c�R���|~����<�7�~����}�[������D��������6~��_�寘E�t��\���k�<w���na��]�����C:�-�M���QT��y^�SscX\�Dvn
��lp����u�-���W_�k7714ڇ����aB�yj%��4F��x�D����2�RyYq+�*6�h-c�UF�����5vrR�]$��ՕXM9��̂uA�A��Q���)_�Dob����bf&
+*Q��I�*���eF��TAKB3[t,��+TB��D�ZA�.qD4='��ja"�#u$e$�ܸ7����{�I0]�rZ��a��Dg6�ȋ�p�	D3tjtzThs�S�]��s��3��w�Ӵ��tj�S����<i�O�	���*(iΐԑu�`d����
+l�UlOK��e��nx�ˬs{*�"�����5�E�sއҲ�ATL4U^2�2y�s�UĀ�긨���oCgZ�x��~�ytnS�s��%�;A�GJH�p�u��&�:� �*��`����v��m�-��Iͭ[Ƌ��g��f�1��&������ ſ�rf�Mժ ��9ť��������"�x>�����
�8q��19e��'`�
���>T��XT���)؛j7G�i��g���]I��J}*�J�1Q�#Aȍ�T�!$Ie��t�WRe&�q`D\4���1}G�2%7���&dF�I��<�k 4�J Ӧ6�1���>§kb]��}��Is�������_o{���u{߂���.~�w~Z��׾���U���x!�9�O�YBI Z�IU���t��Cl=~�Bh��{j�Rz���,m+k�������Gm�����4{^�rlr]��'x���,.+FBRDY��������v�4��f	���˨���l��y-�\�ǅ�("��jKQ��P/�kA62��$��8Di���p�P�zI��eaa�XJn.�/W�����*�^�����P��Loʤ�`5m�:Z�h�GJH�J��CǤ�� %0���W	�#S�p�p�ݦû��.n?�c�t����
��6��V���U����,/�I�j�����<OϏalj#ZO�]�-h�7�u�.��Y�H"���HU��NP�2�F�V��9IG�(]i��0�9�x�����ҷ�dUFg�*r5U��* ��ܴSb���XQI1�k	��&4wkRi�qz=�գ�x��´��,M�P9jLO�m�RnV M���DU���U\r�ǁ*��]��qxB[<k<RB��s�A�lNF,���1$j3�<���zy�w������]=(olFNY9���7"n�L���'Ny���'��Ҕ��l�ƘT�jQ��t_S!\ݥ,���TTZ++e�ߦRUU�|���i����5��z}�Ϛ�
?*$7O8RU92H9�`O�s(����~���&u^ӄ����%��FWWMjn��cpn���A�@�I�N������/��Ջ�Ϻ�oA$�����M|�ۿ������W~����"#���,�x���Jh��h�.Au��>���x`j��.onҖx��������p 6�?L�þ��@k��B5a��o����;4H_VS��+)�i�����PRiu�2�6UA�X�t6��W����Њ�t��|�r�eT7W���N9�9H�KC�QTbB�K\4�/& *!�	�NJD"�PzA���Q���h���XY��#\�e�6G 	@��G��c���4>$��Ȥ�V�o��Q�Hˌ�-)��Ӯ��ĵ[[�q�*nݻN0�����'*��t�76�F5��J%�D�,OP��46�0D(s;Lu:���n���ʳ�íRaT�J��b����4%��q�ӻ�O:!Mt4)�(esڒ�1�%�n�J�'?>��1�y����'hf�o�L<�2��S��T9�i�����H�``R�5����܈��.�L>���af�p�)6���)�Ɔfx�u\eP����q��]�}|Ϙ�K��+5g�p<�y��f��R�x,e�&��!��-�=����!�I�ƨ"�j�"A��u�����k�˨�x��'�R &%I��b��� �C��ԞI�/  �b�N~$4�4��Ջ�,�� #X)Y��`5���פr�5A`h(�����f�ʝ��T"Q�]em%�eML�0c��D����d<nv<�����z���a�#���vlC�����!^S�s��f�047���y��E��݅����_}��~��������������{��o����~��x���:�t��1�WJj��,#��k7����w�����-F>�[䅾2�N��cx��=�P-x������v�^�����z���+�&|�L>�c��'�O�6d]*@zn���^@���JT7բ��M]�f%L-���ӌFB�����V�X����2~fA&/�$Ĥƛ��S��B %�mbF��	�R��mCC��5�
K�O̘��}Vh8z�S̀�fUDs������S�$W=����x氺1K��c��2��A]%�����M��cm��Z���}�*��Y襺���T;������iA�`�{���]��v-�Pb��T�u��S���*h�$E_o��Q�F���1�۶��h��)3VQ��¡��TIy��1%}�Z�H�{J3i\���sTDZP���>M��䢰HKIT��\��ڟk������!��	�!��,�M�q�ekW�	�u\'�o���Q�Z�z��Ml\��1)V���	",����(_�:�J��yNh�Q����9�_)B)3)�����|���ִ��~��t�JȼK�Hdp �h_م �g�<y�/��>�A`�/B�T�!��_�{$�' 9;�X��Ԝ$���ة�9�>1=I�f���� 0a�1f9O*⤤X�w4a�J���1�1fn�Ǚ�˙
괫+�;8��)��E�a�36���1Bh]��XV ��ɕ5v�������3s��"�&�;>���1ӷO�%**y��W�W������}���ǿ����5����?���;�e*��o�����0IG<�i:܉�uLnna�э;X&��>|D�oR}S�J�"�����q��/��4���bϞb�`��C�=�x8�BU6)�_Rs�TV�<5�PUrZ����ꧭ��jG��f-Q�KX�����@z�U5��rC%��J�|�&�f)S3����R�6%;��-+�1i|hr�Ng(�oA$�f �m�K4M�H}jnӴF�sK��4��g�qe	�[���"�blmk��O`v~�=nCO_#:����^���b�W�Q�d<��E���A+�
<Z�!Ps�TڭE��	WX["��c�� ҿ��Ȏ�g����{f���&O�ZO��Z�Z���M˛�I	H�BH�j.�R���D+4�j����r4�U����,��?L(O�D���$���+77�IȬ��0�ZZ_�q�T�kT�+*XPi�4U��ٛ�Aj�
!�S�<�i �ג�F<ޓ����x�[a��^�Ԅ�<#b"M?A����T���������!�B}	���z���G��H*�hĦ�!.-�J_�#��V�E�k�4�Xlr,��"��LK���+�`p9��Wx)�TH*�?�@ᤓ��T~�C}��!8��#����2ոjs� ڇF�������2��!�
���Yh��i�*j]TPJ[�|~p|_{l�q{o��-�����ů~�����2~������������?�����zr���4F�0�odu	��jf�nb��m���9�Clݻke�F043jZ��O�1�\��|����K�^��@}{l^�Q�?u�H}-����I(�������Z��Q�P��rn	!*���F�Ru�3����k��h@c?i�V��at��YE����L^�T@�附a�٦��$#�xD���^S��_DVU$�&e4�8��yUsM�qͷ���(C���Q�>����j��\���
TV8���OGfVR�d�b�"��P�?�4�����W����Z�RV�qk�̧��Dv��H�9՘Ӥ�,U^47*��I��mvAM>/����YD�ajt¥�BL���t�����,�V�ef?ii����>L΍e�4B�VꦉU  ��IDATjx�cO_���Yn5�ˀHpR:U-�,*��s�\�) 2��F�"������2�����R3� �b�_P�!�"���������Q�ᦽ�E����D$���2:�ii<'r.e!� �i�R2�.��'".%�
)����	���Gie%��i��:$0h9G�w�&k�c�����#'�s�>�vsCJn�{�����a�+�]���C8YՐ�L3X��3���F�C�h��3%��˥��7>�������^�~��}�������&>��/�kTE���?�Ҿ������g�vc��˸��9J�9��N(]�a4w�&������X�Eut��lD�f�x�P���7�֛��N�c���˿�Wv~�0ډ������#�-�ʶӲ���Pie	:�:086���.�t6���݃�����]�n���|܎~:��Y� ��׆F*����ȧ�N�����Ĵ���H0J��#��QXY��*�!Fe�V���X�W�F*� �D�s����(A$�h)�V��V��*���	��d�f^DbJcOg����~�(@�@�E'�&��@��l�Z+�L1��nG=��*AB���A�q�w`d��+;n��	�}�M��:�d@�����zګ������Z P�����"����R�)If9���2T�U����M5fݜ��.��T�3����6�flLoE��y@Șc��ϩ�H[=�����,aG��������T'��1�{S'v�W��n ���R2�̈́RMi���T����,/0VX�����V�r�(,c�,GX	Zz�0�/�C{O;z����� _��9��q�����W���ϸ��U�_ڳ�O�Fz~�̨)�n�@}W/z&�{�x�1���})'Y?!$)5'����6K�,T���?�I|��<��|{����o	D_������?���o����|�?}o�m,^eT�qpq#+�TE*ü����F�nb��-\���x���GGxb���cT7�n^���W���W^�^~�ط7v��A�iV̔�	ᅧ+��C��R�1OΏb�
klf �3���atZփ��^O҆~�&��G uH�� K�[�C�dF�(���R����\��B%A�:h�ڏ�mj��.�L�N�H�9�Ȓ�c$>��=܍��FT�iq�B�1�U[$-2����HFáT;���SR+���0:�`�6L�"g�CR$�N�js z@���v�T��"Ϩ��&8��	:��5u��"���0z�Ԭ�,`���@�����w1��w,5�EM=�H�U姹PZkI�?-�,i�t������Lz8�{������3�|�����ʻ��	�]����vaìQ�
,Վ<�<�
NT��@����������&)FJ�i�(�R���mJTOA�i2�RDD�bb�����.���wWh<��*ׯ-EI]��K�QQ�O+@ymߗ�����bPv���J���yz���yAm��D5���q*'�N�l������־~�ON����&%'�3��d�pJ�	H�S�F1�#st��#h4�#�tw��r�O~�3���_���޷ ���w����:>��/:��W������������������_��>���:'��?����M/mb|���4�e��f�7q���޸�ޱq4��ap��ևɩ1��!gd���уع�e�ٻ{m��;��@���ܕ�� :�x:��%F2�-��� f�h#� ��g����bj|��{���F1<5�!�Lꨃ
��Ziu�)���+`�ɋ>+i�f_*F~�eU������z�����m��4{D�%��f��X��i��&��7�E%T���"ӛ/+��-#�D�jkݦh�Uz
2鸲EgIQ*͙�����tc"��B�� ���`��3E�K�ܑm�$�q:{-�-���Ԋ�(� 2�Y����6� ��w��f��Dֿ+�I��3/F�_ -[�m���5���̪����>��M�.�(����D��4����<\*-4
����ʈ��4U���Q�����E��:.dIũ��B�M Z x�<�����阑1հ�s��=�*x��]$1*"��~�q]�H�o��QH��Gj
a�����<�U�^9���h����Xu�e^��hl/C}k�KPQ�*�"��:��At��"2.��<.'���ZbD��q{*���m�s�>|`��C����V�d4����TF#�B�/E$Ii�x��QC*fh%��Ǳ���bgAĠq���������/|��~���D��?�+~�k_���E|쳟��?����]���s|��G����W��˸��CQ���g�0����U�p�NB7�j��뷰y�!�=x��7023�Ɩ&tvw�v4#�t�	���ti�?hC 	B������z_�sphd AAI��
^<��=Xٜ��
���c�K�`�0a�4l�RQ�3�nyt�0�F{o3�k��W\�ȳ���HY��C5Tp�%�uDM}ZwHy�%�V�)ե���j���6�~�,�L02ttF�b��iF�cTqQkG#�+�M�duIxⴄF|�I9�'FB��dt����ܼf�RQ.
/��2���MG��c%*&*��~>�Z2���|ptT�mQ!�S��.3 ���yL�H�y6{�o�n?' ۆ�Ǝ��UY�~s�*d����NJM2eޙZ�[��dt�*n���tlAtј�( ���Rij��L��A�/J�M=UDDR�� �~��m �ی2���Ь�;���惩�`[w;��JS5�ԜH�"㢌:ҘQ���i��PRR�3ӑ_�Iޥ�\[N�s�Z~��i誣��B][��r4�������	Cc�����p���$p�t����qִ:d{y�lO�0E	޽�:��T���}p��kFqM=Z�̘��ӯ"�F���VP�J�*!������g T�Јʦf����{h��_�ƍk���~���m{���u{߂����������֧>��|�-���'����m|��_�o��7�o��Y��wnmTGSs��
�ַ��d�TG�1�qWo]}�W�=dT����Fbh%��	���V��!�ў�[}�C�;w���{w����������RSk�(Fl��At8Ѩ�.��xVǱ�>���)�����QLbb����d�������%Zr�J���R�W���e��nk����֨�~
����oρ�1�观�*nl� �&����(��#���2�����~��CUg�22������J(L��M��IH���W5Ul�)�V��֖Q���:� HJ�(��,�E�ǢX~���A$��YSv����+2�Br3�*\������6�Uޝ���}��L�$��2�t�HM6�vqt�Ѫ�9�m,�ʤ��U��,�T�6�^s?D�?�5�<�i �V����a��Gy�e���wJJO6��$}_"��cL�o�{�Z�n��5V��]-�֜��t4���=�<�[�.BOe�E�O�	�8f��gl�2�X��ҙT(��!��Gaρxe��l+���N4"��M�j�@�L�G2e٦ a֌	F�Ӵ)t���ԝ�Smg��8~��� Suk����i����7�}��� z���-�����_���ⓟ��'�:A��G_���W���5|�7_�}�k_��O������57���qth�Q%����	8����ͫ��a��=�߾O���۷y!n��mCZA.�-��Vs��c���Y���{������]TF{����2c�/x>��
���"�@YE>zx�m�auS�&0>�OGҏ����4l��Dgo�CˢsZg���Ra�eUT�����ͼH:M�\�����I�<�4x���Y��� �%��"53�Ak;�[E���HE��AcV�Bdt0�N�����Zph��������Q{#����J��L���%#b�& Y�f�(+0�5�n{l�%�*���-ۃ�����Ț*�w���2�s̜���P��m�Qf.�V.�4z�'tb�"���\��`3�uZ=4�**��Kuh��
�C�����	��H=�~�����kj��f
��~�*���,]�u^
.�yY�r�ڬW�<��֡���B*� ��l1j�k���H�ӈ^H�':00ڂ��&��sKC���RƠΗ���:Gq����������8|���q[�<`�q;ll`�t�i�FW.7����������!� ��E	�4��$������ߘ�}?K�_^�e��ף����y����]����{��{��oA���=~����'�����x��c�zp�>r��������"�|�5<��k����������N�����w����"��W0�����7Li��L���l޿�m�12���*��VH�hhoBE]R�Sq�����N��v���=��g�.3�t��>�HNj����p9U?:� :�pe0�����0�ק��f1u0����:y��7]FYU9��+Q|�%�TA�Z�S`�P�ގFFf#��, �^�#y>����'!�?�������p2�����	�t����7>�A`�/�B�L
�5���繏��T��t��AD���~A��� �p���"�!�5U˩���o�	����M@T��E�����2��;O�UȠ��|���K��T9��*&� ��Dqy)ꛛ�^��PMOaj�rL�"s��mR�Ϥ㞵���T� �u��eT��_T`:Zg�e�.�1*��T�6+���Զՠ��}#m��&���:���� �W�1>�Be����N����;�o��C����9��N*X�eP��o'��.�;�� ڋ�dPx� \�նu0Pk3J����jg
CsK[\5�7��T�mM��ԑ��68����6� B����V��˗�U65Q�������Σ��o�:��� z���/�~�����}���O�c�����^���������xH ]�w�@����w�p�&�o�oim���Դдu����"�W�0�eQF+�,��0�����|���/Q�� �r��Ī	�嵗�s)���5w��ѣ��Hl��}ط߆۽8p�6�vJ68�p�]����Gx�ƒ��hƑz��6�}`c��Wz����Qa%*��Z\��G��^5-���,���Z�����(!;�/��y)c|�t�3��SA4%�X���@��^P��ɧj
J�x����ͅ����K�
oow��b�^��xi1<�qo��Rk	�LN�:6�,�Lj�9�?��3 ;b1� �K�4[�y����r��J#��H���"oƼ}	�V�����o�j�Q�c����x��/�^�Gz6At���E3�����G�R��ԡ�����c*L�T���mh��A4:9f֘RjP�����:aT��{�ؖL��*����cm1��ztB#Sݘ����b/����]���`��i���@����c<�'�r�����a��2U�66;M�+_���Ç��퍘�$S�T46���-��ռ�elhӚ]���#��X����PS� j:�P��-�rҋJ�]Zf�PQu5�;:0D?��!-G#��o}����o{���u{_������/~'�>��OFo��	�k�vkè��OT���iu���O`��ڧ�Q7ЇzZ��0�&&���71{�f�\ż�4�s��$�>y��{wI��D,BR��~5.�W"5/ݤ ��x�8��c8p���с����`����w`��AF�'���L��0�#K�.�	aHϺh�3�0���6�um=ͨk*3�I�U5� �����[PK�DMTCm���F��P��hp: 99�ZT���s�8'9���; �vV��	��m1���3��2�U�#��>t�Z�G�R��Ϛ�A�ng����{��]��_�@���.��T���!)9��+X �[�p�0�!����>G��.Q-YA)�F����1����dL%�V���c)��k��YOIx�i%W�C�(4:��	TY(�~V#��*��Q�ϪPA �#��Cݻ-A�S3Ǒ�=cs����;���לl��3c@�hzύLN���� j �.�RY	aT�,�H�-9#�J&�R������De�!�0%%�$���G�§p������q�؇�o���6���{y�mq�n?���ue��6/�z���36�ʎ�yA�ۤ㎜8	��H��A1AQp��-�mO��<��[F���L�m ��ʴ{Ƨ�1<�kh�A���j:�M*����@(1'�������S��a|~΀H��;TE����|�����#�������|�s���?�6^�5��ɷ���'���VUto��V�r����1�A֭.̣yh����o֌j���<AG�0�����7�)e��ɯw�c��c�~�M���z��W�4���C^I�)_���~���"���R����C�s�;���8�t��QFz�TI^
@xD��(I�uyIt�]�uo�*�Q�P�QA���J������ކ�v�DtU���i��v,�+���hf����5���ۤ��i�<�>E�r@ktH�Y-��L��&�f��ӘX����$F&�12>���t�t�����X�ʵ�q�
���9o�{zB�c���
�NZ�����ӄ����P�����:���J�����m`XU�����v��Y�<�,���� MZN�
�P�~��\�{�������@8����K��x�ᬏ�y~��
��@L�E�f��D]M��aߏ�	K7�ɹyL�f\�j�ɔ�Ϙ6@�i*e�R�Wg�xmW�x^�!�6�|x.hM��^���L�.aji�Jf�#�o�BE}3�+k�_Z��"$ge#.%��MNEd|�	�,*���2*�>Z:W�w�����'P���#����Q�Q��<~Ǐ��s{q��́}��o���ڻ��;���.�8t��:�����&|��Q�kt`n=�L'!�=�����;C ��g�9����w�=�O?��^T�u������SV���"Ħg!%7Y���6���C���P�;���G��o�����
���>�w�;ѧ?�q|�3�[oD����{�!�n]��$Tf��r�����f����&�yr΢cl�'*;���Oc�0:Ǧ10����L�maj�
f��a����;�=��}���Op�ѫ�⮎'nZQ�

�������I�������)�{���9|Ф�:@03��{m]=N��O3_FKa�z#$ܗ*�UE 2s㨈.1���4!�����:���&¨��Zs���E��cD<�h�NEpad;K(k+�L�-�tX�	�Ñ�#z�����d�K�lqJ�E���N��W����,6���z�o;7O�Ǖ&I�P%p9k:*�w D�Cv���@d ĭ�zN ���!�����c+���� �ڳ�y�Q�ZӃV���V��{Z:@P�=�N=ݞt��ӒTJ�G��~O�C4ϫ���������"�7T�y6S]t���F�� ��G1AE<9Ge�sE �[��֊������������^���9b�%RD|_��s4-�7I�MPq������MM(a`T$�OˡjP۩�L:��h%(��FO3�����]���t���Ö
�f���g�	��ڎ�:9F�~�=����{w�=���������n#�݇�x|N8��9_�%�"�AaMO?�Qt�3��2��n�sr�*@����S��,����D���j�DQM�K+�Z� 3��P����SB��V��I*�U\���P�D����~�cD����ѷ~��&5'�ا��[�x��M<z�Uܸ�jh�4#m���	օ��!cu��40���a���Tut��]@@���yr�Q�Q!��N��T�0{�:6��6�?2`ڸ���[�lkGFI��s����X���ċ�"������#�������:�]{�3��3�DL;�q��N�8���=J(E�GD��%E"#'����g�;k_.����L2����c�X�B��Ԝ����h1�Ac�����(�-Q5�k��uF�����u(��3��"�&'�4�h�0R�B�@7��Qz���i���}N��us'|,��&�@���#�4�BJm��ϻ �m�����@�m�x��Z�m���N��;�觙����YA���LK��;�<���u��g��5!W�N
��� r:� E���""!�㹍e�����*Դ6����T�=�}����(��x\����Ǭ��b�A�A��N�����?W	$Z+T�Ʈan����=��N
:$�i��V���167@މƎ:�U�����V���b��J�tu�I�3`5ARa1��(o�CT5�`�طǆ :����*�&��������q`�+ؽ��x�%�ڵ66{�w���^��{�:uGq��!���..G}�P��	���M�P�tLLD�FI	F��h1cE�}�F	�v����E��H+,��Axb*�R2p1;�@�Re5jZ��3���S�Qw�U\�u7��ƣW����C�Hͽ���w��������6�Ȍ}�m���7�������'f�p���������IJ�@(Uv��rk��I(����Q�x���fY.�t��R��8�g���f6y�^��5*��뷷�����Ul>~��\jjDlN�����œ9�1q�	�۹�p:�A�������'gF̧��H����Y��t���+Bϛ�����>���H�L@y�%t�5����k�غ�����?��"V�l F2�Wu�"�ۅm�}��s��J�Mm��&���	$5�%�F��?ԋ��&T�V�R�%3y12:
��y�\\݌�UсL]���X�W4ݷ.� {��kz��笰2��)�ށ�u~�;
�����,zr�k�l��:2���B>v\�QwW��{.���d�	�H��$:�K�h�cTފ־t��E�&����A�Q�DZGhJ�%�TzMųB�l@#��Y��Ya�"SG��u)'n�T��@����RR����EsGꛫ��U���v��2GN�C.��B���>�*��ىÇl���$�;�CTB�lv���||�vq�Ptv�݃]66س� v�ۏ����v�������H#���y���ZG'Ъkwn�(")�.�*#�@T�7� �u�}�Ե�Ԇ�Z$� ����m6B�@�E$�!%���U��m}�T�s��<&�r�\�}7n��ko��?����� �{���A����>��O���G?I5�����#�p��ܸwǬϯ&GgU�9��v�4֣���֌�����%MU*'�ԁ���4�=mF%5H�/��;�%��[�s�lgoL�c�6�u���Ⱥ\���LD&k��l$e� :!�����3���v� ��+N9��k��tNy��U��(N8��R:w�39o�B#�i폸�P�]JACK9��:��6��7��]����x[�7�v� �\���*m+˄�߿��U��UF��o�6-��p�çfMĭ�2RD��TD}Q�:[P�P���2��� 6!��A�>�^pv9cJ�� :��w�d���O�(�3���� ��;R��|��ͳcI�@�2��<3����l�~���ԣ�:��ᣪ��I;j��1&:8p����g�����^����l䕖��� j'�z;�9����
���1�΍cl��hQ�u�0���3MK�E��SE���Y�P�Ġc�ϯ�yc<?t��_�-�e<��g�ܷ?+�S����H:{k��� �ۅ�{�o���(��Cj|���9���ُ�Gp�6{wR���C�P�GӮ=�	|h�^|h���s��`��8���T2`������1�/�	<]TBfL����������j!]��T?�LFQ9R�*���lDR�DaTDs
�_�����Z*bV˴/�:�gp�N��-���?�6��o���~���D?��?���w��/�">��7���^�ko���o���=6�%k	eE|�t�3�&-W��A 5H�&�oEE[;R�QBEdQE�5�T׈ҦVT3�j�B;Od�5~$I%-P�M���;X|�+a����f��0@9���(+�R?.%�Qm�.�!,:	�	SUO\<�㴫']�`�	G��	"F�J�0��=!�x���8�� O���T�L��'�|	�J��	(*�4�	�v`va�W�ME���4n��\'�VͺA��r0sTH�ѻL���#j��=�2��Z�@�e ���P�����7բ��A�����h> (���������1����:�o dǿ  ��V��~�3rV;�ԟ)�@O�k�nhOǏ���Y!�n3E�������v�;���x7��c?a�H��NS9���޾8����h���+()EE]-�x.��t��Z{hb#3#���� ����A4aҩ�+*`�x,yLg�t�h��3XY��Ma��Yߘ��&���\�¾zcW�Oa��A4���N�^F}c�r�zg\������}/a��a�S��"X�����a�ُ�{m�I�	B�U�`�6{�`��=�C�k/~a�>|h�!�:�c�@-(.�%��20���Ytm[�̒���9���t�*��16i�α)4B�]}���QT߄��zd�V 1����BDr:ᓂ`���#�e�U�TG?�� �{��x�~� �^\����;�p��=|�3�����y������=��?���+_��W�1��?�B�!�=yhf7��Rc!�����)˧'�62�H��j�	��M=O��6��rK*TDSj�����i6'l�TT�m� Z���InRv*f�z�RI7�`��,ܼ������Ul=z�wbbu�A?�.�!:�*�PJH�E|
ᔜ���L��$�BH�B"�H�䙳�#�lN㈝ѱ8|��Q:<g����Y�3��L�~�
DDL"���b���܂dT�����K��n������xm��(�����	/�kE��V���iisJ�i�'�E̍DTC�TC�P��D#[�Pz�Y�HR˗����T}�`���]��D������ӄ��屝��m ��k+hY!`UND�B�`��0�kf9��g�aM�	4A���m(Z՘��M�ު�ޭ���g)�F�PI�C���o�����|^*ɒ�;JlM˩XAE
RC^�����s"�1�<_Ґ����r�h�FMs����5؃�1���hh�Nrf�(�1�My̤����0��4+3>��RKe������\�ƭ;��`w�/�q��gIkKU��:陡g��p��W)�ޗ��	�W`k���ā/���s�A�����ǸG��];�k���J���;w��޽��{�~�xņ�/�:���N��<���l^�m�x/�VQ�0����93��>2I8�'��M�:#L���c��8���Q�ލ2� �%��q������$���6(���PbN!r˫��'�ZF�;6��	U�RBӋX��iRsW��_�U����D?��}�����?����5<$�T5�U�@dRs��`�&�
/�)F�#TE��k�.V��D���f�1�Rz����ֺ�&��
x��W�8)�Rd�>2a
�7�`�0��z���w�t�>V�R�{���O���U��f����1d_��B�E��t��$!"!�TRV>��2��s��p���1�Z:�J�SN.�wt��>��a�p
'�$�\�qVF�=��<��A�䉰���RJ�<���������Lttט�����+�ؼ��o��֍^hTK���-��W]/�Lx���SK����	��:�yMhh��"*DJz�i����\"����{�L�T�J�3��-'i�A!��X@2&0<5˸�̀H�?Dz흹H�#3J�Y�����,�̌k�s,i�gѻ�Ǖ�SZ�ي<���G�Ǫ���
���'O�oh�WWx���y�#0,�		H��BAi1ATeVn�&���;ҋ��A�j]"�-�A��j������籸���k�X�1^���5*�;Vp��,���.��ף��ť	�K��y?�_�}�Ǉ�s���];�
g�1������	������wp�G��ơCRI�w{^�ν���f7v�Ӵ�f�g������^��s'Nz�4.�������8:'�1�����5��k�4����
�h}
!������:^�*B�(�R�I�iH�?O ����dS���T��E�U�뽦�-��.��.��W1���QUҔ}��������^��總�A�#���?�۟x�����1�'p��=l޺���u^�Zc� ���96���T�4M�(n��!��bB�����e-��"*�m0�:+�
k�Mڮ���Q�$�4�!�cR�Lh���w�x����Ǹ��u���`��#,S-�N#��t�_�n0%�J("S�:|�񏊃_D,|B#�y!^���C��u��R19����؞:�c'�=e��?}���ա���#|.(��Fs�b�BT\ "��dQq������pd�_Die��p�3؀ѩN*�!�h�����F��9�խI�nNaae����G�&Q�j���et�i��
�Y��8CE��-�����KuwR��^j��pԞ��ݢb�m$V��Dֲq�"�:O�:F$5t�EED8IY+�, r�����U�W]�p�Lǂ���W�������@�H��1>3���I
sT�sT�sXޜ�ʖ�'�ƕ;sX�9��+�S'S#&�Pۜ���	H�Fd�;���^�4*�ï�I��;�s�����8n{�[�\BTF{����{vbUΞ��+/q��/�݉��bϡ�ܪ�`>�kv�S��g"��ۺ���%.oB]��66��qS~�Du�28b� ���T>����V��0
�2�ªz��K�-DlF�Q;F��%�t�^c*J��B��cRu*�V��J�UQ��މ�����hBs��W����h��5�}x���������=���w����_�G�zbRs�^l��jn��S��r���9�� A��>tvP���Y���zh�M�P���рI�G������
��%���Ue{������3�~� i�
h�
Ie��THZzb��]��y���`��]�����PO���׀it�%g- ���G@d<��x�D&�/$
��8B@����<p�,�t������4O:ѹ��cu�������#\��������m{#8�a�tB����&��d�bJ(Ҳ�QR����*�vV���S�t`j��4��]5�Ȣ���?�iVi-)/@j�Q�"��<j�/9�>.�����=EG�`oT��c[���	:u36fQCr�ώ��"�Yǅԟ�ڧ��a�!���j9[BH�9��K�`A@r?�A0��_��(�ܟyE��\S�֮FO�S�Z��Y������1�HˍP�L�bh��9(�HBf~�}q����o:��A�������9���{����}�m���TAx G��0�����v�<����ٵ� ���ݴ]f��~H�9vڿ�"z��!�8t�N�\�AplrKP�1���YϮbtyC�W0�B-m�wnA�:<����1�֪u@E���링ꧺ���v�/� ��ɹ������4�*�� /2��$���BR�N�8�#ҸPMG���U�R}���T����T�b�n�_��O����}��~���D?���G���Oy�5��	���4�B��|e�����a`n]��C��MphL���H�9���$��b�|lTл,����@�C0�ܪZ�5�L�3j2�v�Y$�V60������X#��n?����X���x�66�J���ʣǦ
�f��(ilAzI9b2s���@^@!qɼ�Rx�&" �pb4��`B)8���p�񁃇;N���ٟ����I؛��#�t�N��B��WOwBɛ�������� ���RJ�`$���D*�$���2UuŨi(Amc)�۫�.ὃ��g^O�YB����u�QTZHu���Px_���s�ptu�qB�As��(����G�Vv�j�ȉcDt�ώ�(�o"��ԡ�ұ��HcE��\��|�:x�VC�FY�u��]�{��B�D��$u��ԧ����_��C����X3�IJ/'"#G�nx�B�ixz����t����y�sv9'�����ۦ4�1*��vTuT>G�ö{����ثq!�ɵ;v�2�s���;w�1-w��j�A��O8�ہ�ߍ����3���LDNEz'	�5L�����mί�ypt��J�F#�W�7����y�/�ux��TCTG�h��D=��£��'����������LD@a��݁�f� ���T�LD<ߛZP�����+e Z��aT�R{R�Ԟ�1S��1���9̭,�j�?��w�~�D?��}"�w�����W>���z����#���3 Z�	LuO2�D}oj:��\"U͕6��D<�	�IY-W�L������sY��Ȫ�Fv_��G	'ةP��8&x!-�]�#���FR��}s��7�~�.6<0PZ�s+TJ��SA��}�ļK���A8�R`\�ig�����4��V��b��B����!��������M�v�ɓNX�X��SNtD�Y:X9[��bq�t������.тHL|�YA419ɩ�f֤�h��-M����B�ԗ�RIᕊ�K٨�.7�t�cT�R���*\�\���l��s"�H���/)':`'�38�"UG�(��`������-Ad���vJN`R�N);��2t��eRu�;����7�5�i���H0-��
���5�ա����˻�N�$"-+��5�q����q:�`�3��	�X�������Ӄ�����+\�:��I{��=j�m�I�!@��`��鼂{_���;����w��;�K*��g����P���ܳo7aKU��e���v�;�q�H+�EQc;j���3;���U��cdu�������/�qhM�S�YD�I�i�A0=�&���u���f\n�gVU -�R�~�h(��xdR@~�1&hf@'1i�,��x���i�')�W��e�(Y�Rs�����R��U�}���oAx�����D:��������؛x��!�������w�vm3��rn� ��W�h��E]w7ew'*�`ʛ[Mz��P�7i7�(�RV��r+,[�.hYƌ,����s�k�]U�l��
,�GU7*�l�A��=��[X���F��1��A�\'|�`��]c�o�p�&��06w��m�0�r�=���)�"/�x^X�IK�ZJH���(x�9>A�O�~�Q�<.��' Ξ���z']<`���%E�4:_�)'g���#�'�I9�i�_�������f���8�)�I���D����e�t?���kY�����MEjv2R2	����Ǆ P���o���̚D>��L+$O7F�g	��bg�R;g5L��rvu6���	�SN��i)Bku�M�N�����ʲ����(��UӶi<K�98ӑ#0�����3�d;��;/_����-A��% µ���g�c	�x�]�IEf.��KZ�E�e&p���L�'��Q|_�k%�0��{~NB(�"B���O��M���Q�j��&��"8̈́RU9Bs�J��!<���u��}�b?A�o{Tp�w^ٷ;�0�o�=r���CG��A�?ƿq���C�����˨j�G��,��V�;�`&����S�L�on}Z��jG	�k�]��Shf׮�!��	�����u[��뵪
9e��(*Bza����e
B�xD'�?B)����5��ZTb�Ҳ����rTT���kyC3�[��d�ݽ&�%�����F�LG����V67p��m��o~��4������v{��{X������_������z�q�&n޽��WL� �*��־�QtD�}&����AT��[��'d^�RnLs��Xvy���9AJꩠ�ь)�H��n�����k2�y�=�C���D��A���5�l��^�N�$���+RL��L�&Uҵ;�ݺ���8��Q���.��!�V��TZ�����4�2NHEdj6"R-���I����q�a����H�������]4~C�B��8}�N�3�ޝ�XR�ؙ��z����>�/�����`DGG"9�`��A���*�q����K��-Fu})j�P�`����Zqy.�2�d�$pZn:qZ㈎;�N<(�����oxS�i)	-+��%\ܜq��ʅ��Ҝ���Y*������y=�H������G�tV����G�:��	f���L������)�?{����̤S� �0 0�����5�?Ғ���Sc��Nhgh��Dd� �09�2�W����l�墨<�(̂�4Sz���d���}A�F�����,<����N�,�g������8����;b��:�%Jv�����C8t�0 D�Q����=6صS����(!s�: 6��9p/:����ƞ�8~��w �����QT׉�>�T/c`f�T��6#K�[Y5�|�(!C��렛N^�>}T|ߠiV:��U�j�y��6��#��꧸��X!�s��ŀ,�*(a��P2O
�{
�P������B�������KH/(An� T�KUՖWQ�F��N��B�h�uc`r�>d� 1�>M��be}�_}���뿖cz�&������D?�l�������?�폾����{�v�:6�m�v6�+T �3�C��%��ۃ��.˲�-m(ilFa=�B�KQ�X@R�c0�}+���uL����������,�20�s�W!X���(o�4a���_���:�661��E�
�*f����5L�_����������},ݸ��-�#��oe�H/�0�	cD*�ŧ8E�� .+1y�5=��b�%���#�j* ,��t��O����yNn�t�j��b"~9mgu�������]���Í�|��Bi£"���*�����T�rM1j�.����=M�hE�`;����ߊN>�j���j�5^&��"���g� �N=>Q�b�O�D!�� $2�l�h,0,�j$����x��2��祸�n���k��< ���,+��ύED<�^b���RsӐY��ܒ\���� �*�P^[���j4vԣ������m�k�E�����(��>��(���P_��{����r���#\]h�pVk�����3�pv����v�S����I1�8e�$��t
��5gI�z�pX���p��*5=���Æ��������'q��)s_��9@���c|���}Du�RX���@��z'0LU3�����et��8��W�%WF��¨yp��~l��h�␩���e3���95H�T���D��Z�7��:w�4�C�O3�	�|�����T� c@��'d *)�i�H�.&�.#��2
+���j�Z��֙%��%����������W�L}�����}�]ݶ_��=���("�?}��|����W���{X�J]]7��&�089���tP5����[0�6���Q��7����(�w c��RsV=5����>CJH��{���X~U���AA����DZ1�Ѡ��F�k]^5f����("AI@2�x����+۝ï[�4ū;���Ѕ,�'gHɢ�s��*���B��������|P(�G#$:�l/�F0����?��y�xz�U�Ń
�ݍ�y�f�.�������Igg8Tz�HUr����әJ��.xt�8�Z�52Q	�����d��˻�I�`�|��|m���㜂4��$!9=�6R�M�+&>�Xt\�b��p*���p1�@�?8�A����PB����!4�r�Td)KFJ:����4*�t����T�g>T2�T~U�.]���W��M˧��+�F&�eҐ�}JCFƆ����Z�U`t#���	8�>	��T3'�>��@�?~��s��S�8jgg�e������R�JI*��������'����Z������	g�;m��\�}���\��?ꢙ���O`ֵ�upC��º�h�s�k|���_°�͢QB-C#�;I3N;��39c�q���:�u���VYs���*�FrA)�M�dQ�i$�b��쓌��#��\`� �h,8F�'UZlj.����Q( U!����C��Һ�m�GEӿ���AM�a� ���*��O��'��D���o
D����?ǧ~�SBRE������-,njb�<��"�T�Ȱ)�l��zQ͓��������HV@Ţ�ۏ��wA�`�BE��!����,`�()˿5cO��ƒT���$U�]V~Z��}����ړ�o�&�/��#hԱaf����+����1kbP���a(�W��k&��{�32L�)4j)j��HUy*o� �vé�T��4$.�T���EÇ��6M9���y! >A!�J��s~�r�Ξ^8��W_�W!�Ψ�������N�	X|����xz^t��T'8��	o��_]�b�󄘞���H��* ��P�i�qxn��2EzN]����J�Z��<?����y�9_3>�	��A����!(������>T�ބ�'��;A{��g���w/�&��۸=��D��͏������qd�/�7����뻶�I����z��:)LfD�9�3@d� 	� @ �@� I�9�0�ɒ,9�,y���lKz~�sN�h8$E���.~V����������CH(�A=3���~�g���������?��=~�������?�W~��_�E�*a��K�,��+����g�4<�/}�s��o�6~����f����m���g�
������	�����������_��|������_��Z��>(�ա���m�ǭ��QC����GΧ���ݸ��M*n��vE[3�:Z�Z�q9��^�� U��!�֕!�����:�������t=!|@
6��G��Z����_YG(���N_����������5�Q�P,!�L i�<��Q1tYrCrB���K+(0��Z4�Yumգ��~����˿)q�g�葧O�����q����g�A��0[;�Q�Ҍ
���M�B�̓X�q$��ň�/D<�(��D+ad���&e���@KZ��M���d�>�0����$9���u�Wd��SQP�d�<��6�1m�cھ������H�H��whĴeҲilK�Ke_4���2�jL���L0�!�>�O���ҟ��/�A�JX�A	Z�f�͐���Wl:���()��^|R}U�z��_4�oXDp�������_�������o㳿�[�U9)�(-��꧜:*O�կSZ�\n����u]Z�����k��9�����>�U�p�%|泿F}����S6�o�1(I�J�Y�L�rf��P��̹_��|�oq�s|]����/s���g��|������'��Rj�����š�����������d����G��*��g��o�Fmv~?��?�_��_¯�����_����{�y}��b���o����(��N�w��/xϿ����?�o��?�g�������s�?��Ǻ�t$�T���M�t�C�<��[P�e �;��2��|�)n�å���6�o��Q��N��nG�>̈́��M���~��+��oEe�A��B�R�>:�d�����K����de�4���?��Q귣?VQ_�s�����C�q �1"Atp��ItBi�L��@(�������\�"��lU5�ں��b;!t��<��Gʐs�D�<}�@�c�_�����]�=�k���Ş�;�cjA�&�����T����!��ĸ�x���q�i�#o�D�G
IL��Ⱥo�8r���~}�<�zF�֣,�8��h]�q�|r�]��T�0�i$�6y���c:��H�*�����8�9���=fYR�VU[�b�r]�M�ȩ�GJab�
y��X�?h�ƥ 06Ŭ�������l�i��J�7�"�Sm�L`	Hj�Ki.8��v�����/���	��ko�/^}�%���3��	������������+-����#��*������ۿ���_�YO7H�)}���į
D�#�8��g�P"�~�3�5��HY���AYs���_2=:��_���/ѡh��_�E#-��:3�#q����&��罖����G\����9����?�g�v�ޟ���yGt8*Z�O*6���)�p�������J��������G����_�_��*��v1���u��/����u���_3�?��3p���x% �	�(�Aic*;���k+j��7��^�5&�ۮ�靖��*��#�M��w�5�\��������zM;�P� �� ��
YU|�*3En�M�����$��Q������l6E��������6��7:��G�������*a�zݒ���FPօF���x�JHHB(�Rx�@���d������NM���,���Zf��2���WQ���jT46���m=ݦ���C��_}�D?�~��	"�����'��|������5���&5�U53p��]����2�V���d:A���2�}Q�29`x"%!FNF����&@i�(o�e�)6Kl�+���0�O���r���o{O-�@Fi5r��ʛ`Z�Q�у��^$��TT�ϧ٭f���.�,X����O�ҦޝZ��P�samr*T�҂��M�T%�S�i������dl�#�b��z#2�h����|�z]KR`T<��-2δ�c�N{5H���U���/R_|����%�[�����W��_x�l��(]���`A��?���?�o�w�e�~��� �������Y���	�_$�>�L�ߑ��~���~�W����|�d��>󛿎���_"0~����
��/�4��/~Fm��y�_�[��?�;���	��J��w36��K��ߩ?��˦��Ͽ��H�D0��f��y�����-��4}��׍�60x��0��9�M$�kl*J���o�����]���e3������| �E���i�S۳�[������Q��-Fu�[QM�S�х��NTvh��ӣ��76��8I��[è�I��}hr���C̚�X���:A��I%�(��O���	D��4Ema�G/@�џ�@�Ś|a��"	�(:�hl����o)���@�o,4.�$&�'�D鄐@���4%)X%Bi�J�.2 J+(4Et�qC�PCg����n�����I�"�D?��ѿ���w���s�0�w7�`�`?�z�=ׅ�f���U����:��ǓBWd�����S��@p�x�������@���W�C�"��!#~��{u.�n���c"�,�ʑV\i\�\��R�e�܏�C�s2j�2n��{���S�d%0Y	d
d:����zc�v��	Y�?������i�+hhBnm�e�)���SpFB��D�)>	�&�1`B�S�'�p�J�H=���bt/z���.8�n� �H����Z �@-���+��j@0�� >!�pΠ͠��t���
�\���k����/���A`�.a��y�FJ���F����?�<�Ǘ^2�C.k�7��/�O��
A�*]�k���_'H�╵�*�c�@����$D��$�ATR*�f�@�k�J@HL<B�0%��%s�F�o�}LLF8��k5n��\�jy�	��&��;փGSo?:����Ksm�>�������j�����S��m2ܤ�.�Lb׋�w�����3�dv�F9.Gj�2O����צ�5)|�F�:�M����/j(n��� �94L�]З�n6hess{�qE�z �5�F/m��{��B��K�%`]D�cl�CvB���DrCʘ�T<�@��`-�o��kZz{���q��-|����Q�F?�~���z$g4{f;��;��۷�1X�ʔ=G�]\���z�T՘?�d�A���<B�@�v'�w"g�#���"g�����-o�xK`Z�ԒT|�vI��JL�T�"�<O�� U�I}wY@	8*�S1�&�p���O�\Jr��ڨ�>뮚���u�N��Dk�� �d-@ը=H;��UY��b�
K+�@"���������4<)�pR��)K�z>�Z>Т���7�_�vHֆN�k�7�
ū�r�?0����B��^[���q|a�z���kL�{m��C3��ß(�Ʀ	r�~�:~�B1 "ڴ���F��<�(�P	#<���	!A5(F@U���G�f���I�!(���و+(B�W��g�*mmG9!R�{�Q��\�C��u�!�˕�v���6B�S�&a@�0%<f=!T�������Euu�Ԡ���lWQvC�vB��h�o�A<2=�	IX��x?^����ưEX�B����J:�C!#�h���"O�I�K���uJRP{�`n������ � ��W�R�_2�!pxCt@�kN2 J�~�	D�NڶD�y&YA0ʯ�jD!T�a�y�{zp������@���3}�A$��w�����Dg�VtF-tFU�|�WvO���:C�CV%���*�R\��¥!!#[LW��-��$G�"����J�Ct:�'eH��zW��wpI�d� ����`��%�g�Sb^�{I�MP|���3=��i|�M�\/$��Z:��Ӈ�-��64S��i�i����Y�VSq]ˠ��#��^��ZO��Lά���"�d^X�4�&��*f<u]��#�U� 7��� c����MXEř�:��uC�SI��y���X��袌� H^�[Q��KtQ_X�'�@�Į@j"��FBME��ڮ��W�#L��[�[�㮏�6��!(�7p=���<�P�0��p9 �](�?��XPv�q�Սt�j��j��4�u���P��Z��5N琢ˤ*�[���p����d��^S�i��Vǧy�ͦՃu-�KK�χ���z�(�]��| K/����GBf�3�P���{J�2ȯ�=W���%�G�^��^���:�h�W�"�u������н�#ҽW� ���k�ib�{.`)}[��~�]�wJg��.�� ���(�T�H7���p~:�h:s���fӷ�����k ��9�Y7Tg��jh��=c����������ӛ> �W������<{ۇvu�5�lFM{���ڄ>�h�^�V��&)�F
�6y�F��`�DjĪ�;_�A���N`�tLAI�!�X0�tGK.�_�)g�)�[:o&��*�%��o+���
H圗s^���z>%�~�+�����RP���*�k:;	�.=[��m����7k`3�>H��f�J��2�����|0�C6�Se�r*�QRKPU!�PûW�����R^�l���Ѽ���K%~H\K�w����u̓��ȧ�@:�Cu�y�#	��\���s�m��um�zt�}�=N���X��[!@u���{WZEبw��4�NFy�����ޢ�6�b§�p.�m���0ŝ����M�U�)MZ�ȣ��u:�g�6��N�+��.W W�h�%Fz-�J�@�<��s�����{�{�,W�f�`���H����oC� �!�	�v^�3������vj��m�mR���>��Q#k�h��;	���|���+A��>rWz������aB�1ڮ�t�z � ���� O I� J7 R������E�&c.���@�� ��o�� ���_~��'�s1?����1���/���"��z�GPi���p��ql؉���Nw��'Ī�f:�&5ԛ���M-��ZP�`Wb���8�b:*��=\0r�zSв���z]X�Ф,�0$#I�k�s�0�)�S �<n�H ��sYۍ�#��Ms�)nT=T,���J���p��J䱓���~V
ߟU� [R��V��*B�� �6�ō�V�z:�S9��U�P.'�'�r�!���{Q�Pq���U!a�W��ŚPXۆ�n�mGA5���ZU���K	��F��f#-���"��PHw�y��M�	�>	�$6��q���ŕ|��[rI5�+���m	�th��enO*�BJi2�r3R��K��D�4yO^5�^%t���f>�X�Bt�%��慂�@�@Huxm��	!5
-jPqZ���!������KiY�>���(-"��P� I���Հ:��TC
B��zD*�w��U��b��6D�a��G8WѨ��5��z�^.%��x���I�7��(���0��pt8t�r�o�������A�5���Bb�i��W�g-��.2�n7��i}MD_� ��D���P�'��	$��(�T<�#:h_GC�k�Hn([�"Ɓ�M�T����ɣ��o�qd	Bޏ��>+&׍��m����&oL���W��p;�v��o3�:���Ո��*�6TR��ǅ��RX:��2>�*+mi�V��#�p:�0=)S��S�\K��Upb�U/�#HO޾
�x�~��ʣ��EH�	^��Y����i=��3��/��������8�0�������^�H�I�qz���i]��Ϧ�y�	f#��Ro�|���=r�* Pr��eUtДq:tWRnM#����/G@�p9�n(���@H�Yj?�`�_%1��r+��뗭gY@&A�JX��i\O'(���KZ�kR��B	DIz�(ѹV#�J�6�*��'� K��������-�ɑҔ)FR��J&���z���^� �!� ��Rj�Yg���J���SJ��b����(�\Xȇ:%d�wGh�`:ki�M��(]Z�F��n�#q{��Ii���Mi�JXN k�|ֆs����	x���0r>�����C�T���7�IIk8%6�j�VEo��z�x�Ӓ6F�n����lݛꈔ��$*���R��fzS�I�"��M��zRPrB^y
�@UHi��&��̣'N�����~��O4}�A�L����������3���V��6��K�u�h���P��`T#�(� J���(� `����#*TE7�Eu�z�\ $�")�@ς��J�!I�F�y�)_ �'p�t�-��o����t�$AL��	�ZO��z��CXey}�/�tTtWa�CM�7��K�'g�Q<]V�\�@�`�D���Σ<7e�>��)'�ٞ���5�
J0i]2��/Iб��Jp�3��%�Jso���[>����zE׺lj�u�]�p�}y^F|���z"�Ɍ��Ā<:^���C7�M�ɇ �_K��%�t��b�͂��� d)��9�(0>��B�o�sK�Ƙ*�hCt�"�
��I�y��Fsd�hn��x�M����V�=� ��f��#�օnܾ�P�|(%%)p9@��"#O��/���`@��De�e���z��"B��)QB'T�Ј*�y�54w�,�A'��?�~:ӧ
D��R���w����at���� j�jB]{�i3P���D����)�uE�z\��4@�}$�$���QHr&��r=D��ad�0�M����$��[B7Tj�d���-�h)P+x�Mh�kwi���D@I�A;AE~t����i�2n9H=����n�`�r�e��H���z g�%�E��I[��݊'M�}��+�G1aG'���v�5G�O:�X�X>xh�֝mf;������s��R[o��ݜ/�_ut��NN�S���q~#�M��T���(��n#L�.[����s?u��=h�s�C�B���ȇ��#� I�$7	 ���\�*b�+D��d�!S��IVp��+�l���y�	����F�i;�#'sNs��M�"�l}XJ^�P��J�	5�h�'��ѹe�߽����?���3�>� �~�_������C���N�)h�z�nAQU-�k�PX- U"�TO����Yl�S�-�M�� �@�VQ�Q�
��G�}݁��f�r�m�\,�|h��K]P,��u�(է�����9h=�s�H���u�TQ�S�QӸL*VS�Zf���Az��f��$�#���uI�r �,��$Z=�'3�0x�u>_ԓ���>F��S`�=�\�A��^E���a���:���9�&:��Q�僄z���
͵�d��9�!a�-8�|�l�!�o*<�nأ�4eS�7�QL�DH��[=�>'�א2{�5�6�((�y���������"� ��d�Gd��^7u=QtAN}����'~U٢8/E%D��U@�u�m]�6d�5�D�#2�C	�tB����2Mq\r��q���_ȇ�
3<LIm����s�0���W��y�����O�4y��$���ˏ�����&��a��6l޾�h�k[�Q��d�Q�:G��"�T�b��J�����tCE���q?&���<�B,������ȼFi=�(����.XF��G�Ҳ]'TwDP�%y��e0�l�2+��nA$�dV�.������GR�V9\־�+��*�:/��"/}&�I���RD)�KE���I&��k�����N�P!�F��m:�60"$	��z�
��'�/Ac���9P2�A��l��R��$�����u�\B�h�}"S��v.{����(�4��R&`b��ˇ�h�����Li=I������HsAHrܜ���kӽ�#"�T4'�
��h5��4VJ�W�|��gq�U;�M��t�Q�"�]uGv�uF����R����"�����I�V���
 �P�6��-+Cy}-�P�ڂ�c������U!$���?}�@�LK?����/�����޹�c���K[��=[�T�a��T�_l`�� O -�q?C-=�[Ex`�<�k٩�	c�#��mcp�䔌[� ʁR<a����2⺤z���-���N��l�����R2����{�uL�:�y��J%�R+F��d+���UZ��b::*��%&��p*BA�b1^�-��Һ��s����a����T��A[߭)�"����m������لx�M�s=)���|���_Et��T�����l��22�<�ɾs�2�ҋy��}���5C)�t�zM߅�/9Y}W@HrE�E��]�\ޢ���FNH"�0 �ȕ��h�t$��z ���l�qw�_iAȂ�B��M�"�M}���F�7
�!�!R�\!��Wӳ��UbB1r�w���R	25�]Kw'Ο�w����q�B��;}*A�i	D?�_��Wq��y��|'O�ctr
�{Gвy3�۔�وR�*אH��*�ω|�+:[���p��XE��O������`�B��ֽ�o�����u����ȉ���>A�&X8���ܒ� ��:%%(9�)���Y�vFNF�7L�6(�Y�W[�f6�,���2:ڮ�=n9tQY�Ȩ�GzU��R<PJ��Eje�Y�d�y���%Z�\��A۝z#��:"���$-+�;E�
�
�R<����2�מ �R��Q�s!l���:�Nꍲ�x�*�S��(�s��t�uI���A���o�(�U+[m���Yc�d��x�ټ�LB9�O�)r>r�a,�:E�` %-%+l�M1YLR�#��rxX��%�8��Enqf����q`�+=��8\���/�4��	B��#�Toݐu5�|������R�HU�Z.��6�Nn�=���|��c����O?���"���D�� �q΀h��i�[�����=2�ޝ;LG�UM*C��0*����WۜBSL�� �^��
s!==B�;��DrH�0}�=�#���\���-�j.w$9sFrK���S����;[NҲ��w�qD��`L�J�TT�O	Ft�����$�9��#�r5� !% e28;@ZZ�crܒ$�y8�4m�<@���5�Z '�!^�'#Ω_Q1�ֵ�

N��K+��[�3)�;�x/�y����[I�VQ�qTs�\]��	��m��-�H�*}[}�媭���+��+/GjFiρ��n�3\�ܜz ��  ���q@I�!��8BG2r��$9��S��&�����uU�"��ϴ �(����'x�Ad��'Q���E�D&'�Wmg�;�3�� ��jǶmܿ������?�Ƕ=TD�[
�Xs����O'�	D?�>��7����8sq��p� ������Q�=���]�����N��Ti}�)��6�Ȧ窍�ӛ���a�@/Y�d��TT'Wf��V��ar�#����A��!9�(�@R��9�[ڮ��Jml��F��JJ�P}��3�l[�l��h�d�;r �F�N{"��B��qkC�)�3I���\0��T|�sHQ�w)�D��J��x�ŀ�d�9�i���@$�8��SҶt:��R^+A�UF���Z+�`�މБ
j	�Z^W��1j1�q@��D��uDD���B���]i;U��������XU}�e>&��$!��x�/|(�� :!h���:�V�jz� �N���-����	 u��b�F$%��!1G}ǩ���EF��+Fqm6m�F��n���������|�����̲T8�&����O�|!���� �	��Oafa�'fqd�9���Q�%�v��C�� ڶlAuKJ=�v�iUE&exT�; �E ������I��e!�p'|��@�\��V�-��6OҢ3�k��ī~E˪or���`v�Ix*�	dgq';�����PrOT�e$w$�$`i]`*�cⲶPz���Ӵ;Z��[�L}���Y-���i��Z�G�2u.���@i[��,x�.��C�eS�E��D�c���u��ӳ�nrC�텡�㎖�$鸩E�t����ىy����ɫMQt�XԀ���Pm�����f��yA�a @,|�GODJ߶��r�r�� ���3��{@�ƂOza�i#��AE5�h����]�رw}|�ܺ{vryߡ���?�o|���*�����S�>} ���D?����U\�y�/���yL����)<<�=�c`�v�	��R_u[w�B���i�0=w���\� v����;��qI�Y9=$��*����O�"ms���#�]su��< rR½_�mql �N�֒(oHI����ɑ�"p	`��)��8u�j������&	��>��$x����#�xQsATץ�p�F�j朿��UϢ���.Gڦ"Yu�Bp�a7*'u��zA��}�vj*i�R�xm�U۸U���5��~G�Cە�Z�-;붸7��@���Tv���|�
����z�Szz ���:'E�)��.(,Q=���\�򷛜+� %/Ǹ���J>8n2}K
>Q{�㊺�w``�0�D'�M���)H�h�L��OOq�ԃ��?� �p��N�`f��DG1q��D�w��;��mE��^�����.��w�is/�7�g�Si�b���z�V�ݒ+�5����A�MnP�� ��uj5�=�^s��l�@��"'��r�T�L�0�us����`�S�����/�͎��)�r�.q��{2��T���t.�1x�0�t�IJ��9�6��[�,-j��C���^W�=o�ɐ�9�k����p���^��Ht+��*.s�>�2:��B�.p��y���9.�>�x�1�;���A��t���p�)�ܬ��7��k�/2�䞴�e@"�|��^@m����s�d�b8:?� AH J�K�=L�=O/,@ny)���p/�=����[Q�ԈڶV�m݂���|���{pra���@dk�lʂ�~�%<��S�>]uD�9 ����7�!A4G7t�'�0y�Ʀ�0>u�F`���Bid����EW�܌��nt����`j4@jEQ]���<���,�h%InA�u9(�NÄ3���(�A�WNvar+����Mʶ��?�#��xy|m_�pes.����N�nɾf_�kF\W�G���(hL*ʳ�K��N���%���emz�vY�"�T%�*	ܦN\�3W�r ���E�c6J�6��ܮ�/�Zt�5{_��#	�e]o�I(���kQ�׵��*3�&�p�k�Ã�z`�,�t_�]�x�\V���4??2�˒����ߩ���� �B�a�I����M�^��x�"�Wn�� dd3��d@D�X.�R"���4\D���t$-k�����YG���ϰ�ƩΘN�4*%ݤe'�^����A��h�Ǧ�N��M(����(��ByC��7ܾ����Ğ��1;���V�Ҕ2�
&p���<}j@��'���ݏ�?��߾���0�8����!tb
c�G�� ���֝��޻��ѦF��{��CeK+6�nA۶�ԳU��(�@{UF�*Hsu��'�8��e�)6�4��&1�1I&X2ɥȱDA*Q8���Ƨ�R�\G�L9�G�������8'�A)��*��6���R���U$�DٶQ������·���f��vR�R�=����K��u79�i���t��[�n�K����B�v7��+�m��[�j
���ԠW��b�
!�B�;�$�7�c�F���'�"	��8B'�	+�'BG
�KDTR2"����S���x���yRV���J�Q�چ6��6wwpy
*J���I@塨��uՄT&�Ѿe3�����]�G������m�㟞���C@4:5�}c#�0?ކ�{>q����#[i�%%�h���u�݄�V4o�C=�K5�Lu�����ɄQR^�i�a��@m ]��+`j��] D��'�r����TAd���w�nj<��\�R$��RNC�մt�,ĝu_=+�}��n�KJ 1�qB�í��s���ђ� $�%|�u�� �@��00>�K�0	!jD�X%s9��!3��9H��Q^Y9���v�ot>�e�H��FbV:Rr��2��� �$��0پ�[�� zA&?��C���;:�������cK;�PKk_��@�SkQ~�2#���t�ZT�@���:��j�:-�+�� �q_٩�&�A��N�,Ff]O�*JR�#Tt�A�@�!+W�<LOD���+(;@ҵ: qzt���B�M��.8��l�9�jac� GOD���}嶿�����c�/|���@�z����҈�nZ����1R�z�H�	�NLA��Q� |\���6���b���L&Y��)��FU�&B���KG$HE&& 6-�8�̢|n/2`*��DY}�S����ck/��ډ]|����O~=D��aϡ�� ��wSW;]Q��ͭ�4ʫ�Bzq��ⷔ�"S'��44��";IPʣCR�u�E��^�wZ�;���f�2]����(�*�m���)�ȑ�7��-@Y�#���C+��m5-�����%�<=�|!�|nߩ��"%��F���*��^G�D@FA�r���4�%+.����-�O�I]=]M���*'�I)V"������2
r��7�;��0��׋��~� �D��h��Eu�ǻ���M��hNn(��܀H�H�R������و��2�qrK��iW��l>S���:�(�a$F��<�t�e���	Hnr���z� r2�$o	D�28������ed!�^��u,m���/&�9r�.W�3��#R��J�&�*�.'��&��	%x�0�G
'|"	���L��o&N�����TWR]k�
�r~y"�	��(���'$�$ť�"9;�H�s�U*��1R�Pus#��m[�� ڽo��`���KW籰��?N���z@���i�@7i��Z㈲�w�`2�"9"�%*�7G���&A!�J��R�Pvy
M�kjM/ �A�������R�ὕmFwd������rY�� �Y�R�Zo�5��1�M
�+��L�>�W�xI˞ �X�D�T��TL'-m_��.��9{�����".�6_�5�}ξ����s}��^��G�����8��^^���	6�V> r�(�"�1g�!�d��I�����%)� >eI��M�^���BVar2P�OTZ����[:�42r.�# ��d���Sg����8���`�bRR�#�T,�]\���R����4 �q@Է}�hn��ۅS�g�O��;6&�A��'?�~�=����t�Ο��iL��\�����Ys�#RFNզF�#wQ]�)����"�q@D�{@$�i/�I.IR�R���R�[�ᤫ���-)��i�A* �� `��>�Tl��-�tliے��O`�ъ��m{�R
�� �%���e�[.+����Q��JX-9o9`yrwP�l���z��^x�o��WZ�^�x���N�߱�|��/ܤ�O�Q�R=�Tܦ���b�Ei]En��. >r?���>�ি!��Pz�K+($Xҍ�	��A@D$����
�D`Qt�qG�PB�Qf:��R=0R��眢���MDm[6���;�vbx� .\<���?ۘ��3�� zR5
D�އOk�|��a �ͰEt1��N�4O���G�r�(E��j�i��^��HV��2�J$����\�<:;�H���0~Fh�g��!�W�[�w��L���L�/��(r��vNV��K q����@�>� Z�������P�)tj40m���: H���+�-/�ΧY%�Oi29O+,��K"	��� Bg]H(���a�AE�"9Ip�+Rjw\j:��i�S,��,�(���#A�g� ._>����٘��3�� zU77-�o����[E
� �S���|���pU��Pm�Tda�&�0��"1�tPK��TTj:W5]�WT#��)M`��Ăběn�	&~��A�����{��܃�{@V0v��S�+����X�;�����r����9�]���{͎>) ҈����U`��nS�A�!���hH��״·�(=�������(���HˉOl:�!|B��@Ȭ�Z�g���B�	"ɮo�@h�-�S����Զȶ)�@JN�r�]\���V�}�q��E��`c�D�|��I@Բ�tR��`��T�SG�"��
%�z`��p.��s�a'$�uch��$�L=�)�$z)tNR�$B+���}b��&� �;��>�z8���X*gc�@��._ 9r���$��]��� G�iP<7i�VoDu��ߨ~��MG����H�PSт�~�9y�]�fd�h� uNg���`Y�5!!x=(������8N�1"���9HR��@�"<9���L�1g@TB�)aAuDn �'���p���A���1�A� �imFe�&�z��j�	�0�8"@N���#�h=�O�Z�c�1:��C�)DV��U7AMlN�qDD��Q�� }�o��դ����v|i��<mw�;�܎aeaaA�+��x�|��"�8��}�a�H�F,�z��Qv(I,N������vAI�
'|TԶ1"�	�u�͚�`���\���	�
5��w��+��o�:!��P�R���q���L7��!����R�
%�{� �}纍~=����/�����р(O�ŔWzR��T�N��(��D��тEg�ʧF�%)�UEtJmV1����=6aqY�U�1N]�'p=8�@K�13�) '��Y�ҥU��R��n��pv5��;_)!�7�ϑ^s�����R�nn�k�o�AK2�+�?�� $�AH��P���}0�q����T��&A�U�|ӗ�"� ��0 2}�q�@�m� ZEʚs���˥�}���"Ӳ����E��t����8e�it�h��W�l|w4���7�~ۛ�M�*�I�=cT�QE�ګv	*U+�(j�nkT���j�VZ[Ů�U�����7��<圜���u����}����ې.�F�D�@U08�yz�,a9���yb��g>Ԝ�)Uڤ1o��������D����������-D�]Iq6�H#0J1վ�����w�U� ���d9��$,N��w=ҶE%����`��e����'��|������w�pueB�&����u���d>��~�iTj �(�
��)�����g%������2�K���SZ��{]c��k�?i&5���X��*�7��12(��?$I땟9,l�Hܟ$v�6�~9���L�-�^�X矌�u����,�\�?�Ć������w��^�����L��g��3���\	�����#�i�˪ҝc��O�D��{J[�Uo$�iz�MuU���k��rؚ)�~�=l���фz���͍�f���y�����AQ#�?�u���x�^��ג7;q����T��T������x���5�X�%����Ǔ!��(��3��~�8�����阭�r:�=nq��5s�ͅ׺�r"�R��n�p��.&ȝ!���k}D�Yz˦�ɲ�8� Ϝʽ���*0�Vf���xǐnXq����wY(tPL��?�q�j�-�.� *l�Ä́(�H��Xv�|��c�u%���#��7lwfGB�}B5n)�����5;C\פQE��d������SO�����e<������R5�����~�t��os�J_��W"14��5U�3��qI��:$O����Wl|��oe74>�ܸJP%)�������T���ť�4�{r��iE8jH���vr|�{v�8��tB���EhS_�iF�M�yɂ�.�V*�F_�]%E�cPDG�b8�!ﲟ�� ���
�O���Z�Bg����e�<����k�zl�����BeD�מ�!����?"óԼ�V%|��DdVQ��[\9LN&p�,�r��G��]�`���_
��*��#D�hl.��<\�!.�������]nV���J&�o�WqyR��ց�J]��݈��Ql���~0��n@�0ޥ����MY��Lq��{?�V:�V"g� 1.vS�Ւ�Y-$���՛���r+q��h�?������K�V؉��}-K�q�H}C�1�P�.��I =�qP�dYo�(�x��k�T���4 j�H�3W�i�{]5�v{Ԙ�c!��������?_3(�	�h�15ØGEC;A� X��Ybpȋ򷽤�2�#j�n�jWS�zct� 2^bW\g�z;�$ ����G���s��-�M�%�C3�51J[-�J��'��¶ɖP��!k�is?KB��C��7n>���ষ}Y���Y{�^�K�����z��;q����{�w��okn0x��S�k�����9��W�W7���O�.J��Ph4*�h�����ֺyR����	B�2�i~������E�^��fV�,�������FǙDRr��מ7�����o�fYڻp���"����E��eRw��ʛ��e�e�{���3~�4�>z�ڔ�Sp����;�3$	��pt�Çĺ:������Nr|:��k\J���Z�&:R�g&����:��;d�A~�'��%�BW�9���a;�w������TOλ�)Й�n(t�~Tl�A�d���u|<5��RdX������hbS��̠�(����5������^��~��p!:���� G
E4*� ��%��(-����"@C��kws�[g�X搴�.��ui�*VS��b��aÑ�o6>�c%�:�[��Ķ-)�����4��ik5���O��܆g� �v���cblUd���_����nW������tN��-�ix��ʆbʏ�!�'}W�����e���_ؠAE���;=��)��Y˟�>��E�ӈ->��5�R��_��e�P�>K5�8��hR��m���OE@�4�t����ŀ�^�F�a!�+^��`��/�(Qr�����9̊l7��k���0׆����
|T0[�_���&	6G*���i�󵭍��k����&�,-*( t�i�=����d��s1�[!�tP�&8���P���ڇR�7
�{��a*�'l����� 7^��z��<;>EWt�3[���jWŃ�d�d��G�?l��V%ޡI��qu=f�����#9��.�`t"�7O�jt����L�5�9��|�v̏�8���qX��u�O8b'�Q�Ո������t,k��N�މ��nu�pO�;%u�rc�MI�u�5��Se�E��ا����;6����p<��?���B#�Oӹ��K��gV��XX��G�q�Ƒ���+_�|X���ʣ6�4�6a��º��C1�]��q�=4`�� ��Û�WK����<�">"�]n�vi5����pʯ�U_�X�c���'�\X�uu�.��k}3n~�,�CBg��|jl<i}�ksq�	.qB�s����W��`�������a�%�Q}&��[*��JR�Kn~� ���IM�)r%;C�o���c�M���ʝ���ժ�(����Q&�+�3��Νξ-�7<
��wu�Ͱ:DR��9�r�q9 
6�$�����۪wЈ�ڟ+3(<��o�S*G���ٽ:l��JRT�V�)��߆�ҥ��]�dj��AK����ߎ��Z^�"�!�$��.��+�
/��&E�a�؄��`��}qG�I-^,{��	x?�' �+���Ce�t:���B�?]𹅩ܻ�S{Q˻���B�e��㱈˙+U�`3�H�؟ugӍ�c2#C!D�K�{�ӆ�c~ƨ&����ls��H�݊�N8w��U��:�@�&*5Z�J��r�'s�q������0���$Ϗ�*%��R�pYf)��%0�� y�5
�)[}Gϥ��w U��E�C���!�N}w�扸�C�r.���!v|��G���;]i��k���0�r��I`.*B$E��~�k޽��*]U��8� ��C����D����ځx~]�Z�w1�g���g�6��̮��.i�ӞoG~�R�W�\P|���]G���:�L�➴���ԆWJa1Tzl�j&�ʅ�Q��Q��Ƃ;�{]���ꙏQ���v��h2�㾵���,��&���� :B�.���&I�u�`���K��J~���{Z	A_r�5��**����\כB�`kĘ��T�g�>DO�� �xNX�|�Zz�j���lv�i�n3-�K��bB����I�m3�%�<�-�!��vN���Fjc���3zK�Z�'k�sՍ�ld��(�M�JD=����ç�f
+��O�%E���D����%kV����Չ�4�|,��O��$gB��3nP$ѳ`�8t�:M\Hjf�'�n� U��g���"�s�2&�~�*�dՕj�Vzq6Q�ξ�$�&b�u��m�l�]7��yn�*'�]����<gh|���6D�,D�=p���k8����PTY4�F�䑦�ܭ�'�6dV��E�s���,��=~+�E���[�<���5��"m���	��DHk�Pls�Kj�kN�D��|֍�~?��'7�ŁqF�8�A�h0S)�s��x=��l'�B껄w��_�~
�ܪ|HY�����xw��d(|L]��3�8��- v�*<�#^�rř���a+7a ��3�@�}�aRұ�)&�����i��3����;+�<�vI��R��n�cP�R�8o&���t�p�T��w_�	����i��l���gB�n��/�}
:~�_q��G�����s��}1z�ӆ�'7�?�f�M�#�H[+����g���q/3���;ܪRY�B��?�V���O�b������,\���'rjo�CH$���0I\�!��vZ�7X���B��В�b��M�.Q�4��E��z�s҃��P%T��w��K���!�+�I�A;N-?P5�� ��zw�h�%�յpX�}�s�_Lԩ�a����J���9�L�ȵw�W��Tn"��x��9����)x\�I��U~T�d��y^'���x2���ҕ�`�G�}
��-Q	]��B���$?���)T-A�@��fE�@��@���2mnG�n�M����Mx�^�fO�����m�G��̏XN�VVzݛ:��~(�e9�;��r��f�ηI2qԵؖEao��4��F%���v7�\�����34�*�K�O�j�����F�E�`�<c;�Mq��Ǥ���,C��־.&��ʣG�_ןyzpu�:Oʫ��+��՟��̤����9�l��}�8�8$�Š�gZ%F� 22�|��Vs��l�Oy�ɦ&�����V
��Q��m_�ԑ�I�Q�&t�.���#��ۼwK��s�H��-�&ڥ ���Û
%M���ȧVU%�(Z���ɣR�R1�����FH<���JesQ0-��;����.��ܡO����Y�I�H$�T�rK����O.�<����a,�tp����� \TeO����|zAZ,�YdmO;������Y��SE9�>KH��ɮ�#���?;�So�ă�iv�8��)^��jAܷ�(0�o��n�sa�]IaK��L��-g��*�k����NG�_����f��=�;F�����j�����{@m�5�@M�� �{~�+}��X}=ۿ�[C%�Uf~��u��2�E@��W���jਟeM"����,��ׂ���)����gm���a��h��0-�w9��}t8VGª�s����L]|�¾٣�w�|�DB�� "��������'���<ҍ'� DRz�	gzޟn+�v꼀)�Y����J5�t�Z�n?47$��w�����o�(W��e���t���O7|�$PZ��-b��E�I44q?�`N"./_���:��.-tX��A
�쏩׽'��2�َ/���)�IX�i�/��A��i֦Ю~����Ae�!y���"���B�G�3���^Q�WD9��Kߧ�?M?��~B�D}1)��O�����4�)�4�Ϛ��Z��L�_��[qD�t�L���ϴ�jZ�����WC~�q��PZ�J-,��d5ނ�> *��X��sc[�n�C:�{{��j��_�����S����D�����^s��E�'vs�-`����9�ÈK3s�����y$����BA�Ƭ��J-|b�Ć�w��AX���M������P���FOٛe+�W�Q!��\�$4Vӹ ��77����F��E���G+k�g'ʗF�Ĥ��zTVɥU���s:�]�9����u%��T�fo�uUQ�2�HRk�1\=�W�&�|w�Kb<z[$R�-U��eG?���� c��h��D���DCh4�yr�U�'�)o�>
.k��ͦ��$(c=
JnbV,�����0��f��x������n�p����:�{��7����+���3w.�`�����J������T�	7~̶J7����-�y��f иd̞�N݉!0$BW���}~��_7�s_��D,1�Y��{+i���;����ѕ{�4>�����*!�U~������27^T�D��:���ۏ�v��c�-xt�)�!_p�T�����C�s,�4|�>��@-=c�'��5w�߸",�իc���7od�~,׶� uت���)�3Tj�"c���0/�K����Ȉ��1�;B�
��?PS�/ȑ_���h	qON8�����ѐZHk����G���vE<
P� �&� �y�n0.B	��7}�c�l��4�����(�U�`�T��W~bݑ���g����o��f��cA�ӷ�����_��ԛ�Ǥ����<e� 9�_籖�	R,gH��u蠔�-OMB?V>C����{(&�gE_\NP�17��E�}��s�\�8:y��YŰ���R�L���%LF�������}���5����o���u�u��y �o���Ҭ. ��PKM�/Ob7��	�����\���+{�{��NaߢN��'0���1!d�N��c�)#�k@3!W����̡\��n�7Z�D2G�~�?�b�� �RYT����������Յ�X{�tv/��4K(^������z� �7�1�`)��>�����lXzC����xy���p�	ms�pS�g�J'NW����2Ċ����\��I��h<�]���H�����nN���Z�p��3����32��?�q.P����]!|�rV��ZW������g�O�2)N�@:]��jt�_���z����u���B�dJف�|���� �	n��
h1j�ͽ�!����O���])���Oo���-�a�7�Ky����<���z�4����q���a�ΓE�_Sǝ���nj�,
95$��<�q�m���T�i�y������oy�!zZA)�h�u.A�˕V$�][�O��`��O�(78����0�|Q[�D�ʼ��$��|t዁�����HQ,��[7� ��-�Zk]n�S������B��\ޣ�d��G\�@��*���U;۷*	go����O�*��H#�n�N�R�w �Fq"��/��
������#�筁�f�`�YI0�� ���1���H6-F�S�3Ĳ��À���c;M4�$�k�L�oUΧ�QX,�(o������D<����ّ��L�*`訤��<_ԩS��Zf��<jm��)@c�$�����$bMA��{��sc�^	s�Z��l���"ƒ�V/��+�v�h�GP.�Ǆ�$��c&(p�h��)"���ͺRpb;z�M��C�X����<ƈ[�m>��sB��i������k��_��(::���n��D6�����>��7'G��kJ�AA��:��ڻ/-_��Z� ��c��'`����H��:A 4�yy���-@�����x�dO��5z�q��&$0�b]+��T#��a@@�����ԩbc�$F��Kp���E�rl5��$���M7D�m���k����1�'=��"	P�9�v눬�x�U�W��I�W��X��.!�V�'���W)�!��4��F�GZ�E�����O<��p$A9u�mbdg��F�9n,��.�����yM���$$��j���v��n�.�ǥ�7}� �U�����~�"Vs�9��Ŕ�/ ���N�Ϸ1���G�/�G�����and(@����aPblb@Wצ!�g�����Y�Lّ�!�b�O4�B�n�RR��V쉳Y�C٘����d�<[�Mz!V��:&bM�2��lC����S��-��B��14��ŚJ\�����5�%��H$������AW�L1@�Ԁ9f������7�dAE}d(;��;��ٸƽ�_�?o=���y����t��vX~��W���kJ�;0"g׹���b�4I����% ����j��i�f�q���,��3=�6�,)�Z�9.�!
��2��] ޼P,�tN� 
����+ae@���"/ȗ���?^�cdc�V�����/���HX9�i�#��������T����/�9 ���;aj�1+<��!)��l2�" �����=���B�,ՈP�y��Aq,�HQGD�p(�!T8�9f�}h7@�)��Ŀ�.�ϟ^�	�`W�y�����.�^�eׂsy/~&Mg���n�S���8���D���|\�W��7!�)ܽ�Wɐ�`�E�¦ f�g�ۊ�!hS���t��t��g.����Q_9E(:m������|00d�k"\��xe����8�%V�O�����(_�M��T|�4�\k�y(WݪW�,�QxS����騤X������?��e�h�ֶE2 2�oi'�y������
:�^=J)����~6B��N�Rz��J�8Y�7���B��{��������fʅOm�}�����ٚ����\�Ay���>2�a2�Wu�g�<�&��i#
=c���pt[�E؇Vc��^z����f>;�	|�ۿ<�O�s����ogo�N�����rF�c��*����H
�^w9���]D���UQD�����x��?�/#2�OK��@Ğ�o�Vh�;��ۿ�c�uhMyt��x�e�6����/�5�y� ��k�+���2Dg��t�s^��v�A����]V��>�k1|��i��2lT�������t�/[(UL-6/��=�����TX�F��+A�+!���(fN����ia�#�0Уz~�G&�P��9���Οe��χ�����٢�b0������Hn�r�Gi ���3���jg�<� ��ˋ�Vz�x��COW���@z�����UA*L�b*Z��ރ�	^��y��G>@Pm/���.�E��]Ʀ���O�11	Fن�|��X]�Npu+�{6����st����o�מĺ�Χv�S^v[4�hTV��
�IO�O�ߨ����v��2�a�K���]P ������F��_ 觃�swSd^�Ź_�>!">�0"ɴݟ� k0Qa��;w��T�^ɸ&�*�oE<�vst��m��!��!��]G�;y�� �T�dxy�arLM�R�8�"o^�m	�Q�����[�H�y��~�����_�_����|^t^M)�7g[��W`�m�io���\�!����Be�T��s3X����� j������\�wWb��`!c`�-��!�YY���*Kv�%����t��	�9`��e�ħ���=�d�f�`ID�<��".o��E������h�1�i�W�q�H�]s5^I��x�"x��Nϴ�?�����A�[�b�lP� ��,�|���cO�.0(R�X9�3M#�zyU�%�S=���%�BCw�H�k��v�����G�_i7ROB���z�+���Hh�Ů��P�Wh�va?e=zJP�e}��t����`�j�G�X�L�9�`M���6�"Ы�����'�(����F$$�<�q�9��Ӹ�oH�#�>�|N���J���U���Leǈ�棱�2^>�@J߰�iӂ7���S|K�l����W�?�^c��.����H��t������p�}���I�D������e���Pμ�J0��g��� ���g(�s��H��R��\^D�H'o�0�wSH�ٯ�cG[�%��9��y��O�.�Ͳ XP�M��Lޯg���$��=Г��D��*��}h+]����Wr�֠��m$�����.�:q>�3z�W>���Jk
ǻ��l
�bA<T0U��	����i{��6y�5��<���7��=�@�1����4�Yo)*JKa� ,��^�@=1-��f��a�!�c0�N�qܯF��c�z|����E+;���;fA^K�����X�9�ܪ���>PP������Fy�9:�2X��7M&a�,���`��9��"�=}�@��A�K:6�X ��y�˰T+���A�h��ez���o׵�~R������Bm{Q%%/|O�`��pn^��&�o�_�I2�� ~���x�ίFqB%
��\7�e�;s�e�WӍ΋�☊?��[~��y:݈��6,"�-T���o0��p����{��rr2冚��&��F����n`V){��\�0{B�� v$�@�f�mo��E��+�64�D�'��[���Ϫg�y��3%���_�]�~%�۵�MQ�������ެ���@5T7H��y댎�Q�s��'�o1�z�.����PIQ����ޠ��	U..`�,/=��/�|GY
�$�&D��%�e�z��U6v�M�q*�d�>A��@e��nr��^%�-IFY��v�0!2߽����b0߰`@Z�U�)�zSn��^�s_�����u����~�1H�ә&XQ�@���ԏu��m��z����m�E���G\XX����-��*�^iF�zㇼE�x����g~���w<�Z�_�Z܌'�G�[_Z`���ܪ���U='�1e1�k^מjj*l�ښ��� �M*'����Ad�*o���3��G'(C��ΟS`Z.�niD��{O^����bn��1�Z�(Q��Y��W��|�Va:v���_"N��t|0M����f�%������M;Q�f�9���O^-���CvH�(W�ǠH��}��{cң�G]�K��JC����g�3&s��|y�Bc!��<|9�i�_��:�p^���O"(/��{��_���|W� ń*P¼���ur��ÍMgΐ��w��(�-�R�����'@0��O����ܖ��*ֹ���e{s��߷-	��_8�G%۝2�}Ni�oj"�a)⠳=�n��j\l�q�f����	��,�ݖ]ɾ`|��52>�\Ï�1��j�ٕ�
 Ε'(���BUڥ�^0�rR>�XZ$������"��(�o��>y:"��%r<���ˀl�k�Aaa���EMr�>t��<���O��.'�+�7�"�U%`ʡ�l+ό46Tٱ���d+䵵�69"�z���0��;�L�7���"�Ox����k_�Yl �m�QK�T���H��pf���;p�rY���J�Q��_!bK;�Z������#��^#��عv짚��d����Gĩ���:V@O9��$M�����!˔��7����)3�+�,�D^��(T�U������D��y��7�V�@�T]]dZ,{��A
R���*�Z��W��7N���r�ə��@�_�k�<�N�=G=w�Û+O!�i)�S�����QǣX�]L�yP�;�{\�S铌S�@�%�h�G(ñ~�7_�{��A��cɵ٩k��0�$y>@�� A�a۪�]�In��IJ�y����4l��T	���Mi(������7��Ms7��n<�+����::��&�8�9a�R�0h��n����]��0wn�_D�]z��4}�>�>y4�x�(��wAdx:# �엧��^�����fG�X�����W�b�hPkQ,t{�d\�����o-!��sދA#��/��-7��X7��F^e@B'�q���Ƭ};�O��ضxº�n��x��q��We|��q'$��b�1S��̌$�PÏ`ܽ�ѯ�@��F�w2�d*�������:9�Z��oT���
Z>-�����Us��E�
C����)�.ۄ���)q��~su�0
A@*��涉��i0:��T�u�����D�w��p�`n��E�ń&���;~��54�B"!�FB6��K�����F5V
ˤ��WD�{g������d����3��|z��j��9���c*��_�p��:��S:���o�����ޘ�S��w��c�0s�N�҆	��s�X#w��wY��Lj�cq{;��b�B�k�k;0�l�����^{Kh/Me<Ik�&��K�u뒶��f��B������'����V#�<���b���J��~d ڥ=Bc�5^�⒤f72E�R2A
d�oH6�����)�a���T�f�*�3p�h��۞p�HC��{ ���;?F5�]����,��L���_8�(
/�>}h��aV� �}�څXS���x����ѡ+	�rǑ�� ���kt�li���~��r�}�T�G���ԃ��D�U
�|�挤Pc�5�w��N\�cdT�t~���`� A\�\�k�3W��]��~��_|���x���N�Ө�	�7�]LN�9�`%̭S_��3�Ɗ4áb����ct���42�����%�7�+�w�q����Z��|8H�K|)3�� /'{�	�&�T}jg�.b r��&]��ꓮ�α���V��;H��Ho�H����e^a�I0��6>��yc���`p!��һr�4�*���w�_��	�כ�^9�æG2����	�1��g�W����'YȺ",���38�e)%L�9�/��>n��<�?"�&���\�����b-!�,?� )3*МS��m`���@����0b@�5O��^ߩ�~O)`5��X��2߁��i�HV>��n�,&�>�D3��N��B;��[OYU�o#����M�}�4�W\;\�V36?�Ps���$���1aR$�Z�"�卡8�d�~5��:��î;�>�$�����BO��A��dF��+yOW��I65?J��޴���8t��O�;b����d����(���GՕ�e��F=�E5������T�K?d
����5�&�9�d�/�r�sp&?�'C��5��O���-�Z([!���7�4a��JK� S';�Cm��H9�Ssv�EG~\�����zDN0�t$��̽���-��f|�v������:��Z#�س� ��mXu�1�G�����ޣt�G�9`�&�ƥk��K�-����b7'�����f~�����Q�hƛK1��X~���Q����Ƥ9F�$�Y��D�Ǯ�������C{,wB�T,f�������������W���In�����T0lx-Ev�k>!��R������3MU3��K]c
�����4Sx�	Ҋ������Q�AI'F�͉ҏyJ��}}W��d2���>�>��r�O��)�#Bi��()���/<C��~��h��3�*��y����D�����r_�Fc�^���ǎ���ͩݜ���O��h���W��]GQ$��c�Ћ�'�y������	#��>W���|J�$�����Gy��J��p�%h�mߣ���'����x\���n�|�FTQ�zW>*�N��o}q���P���dL��F��U,���a��L9�J%�̘	\��]R>r$��-�N_()��! C
3M��fúFL�w������PD�l�P	�8(e�{Hqm���5B�ކg.f�S[_����7�Qt�M��aK<B���3xe�;C��~=�͹%!L�Hn>�PJ����7u���N�4�FQl�72��4��~���<LJ��R�~�$��V�4p�[���?s,�ܟ����x��^T�9�b߇�!�5��Iy
)I\�IF=�-i�~mu��Rӑ��v#��Rk��i)uSS��ݹ�f�q�]�x�k��LRW����ٹ�w�<6�GW��x�(�P������2Ns���gMK]��?�Ddj�>�=�,�'���J��t����M^1�ϗ5�oO���k+�M��_���4�7�����V)C�J<1%N�O:��-�x.��}��e���ϭn<�xQ�cв4��!��������u.�ؔ�G�p����B��D��(�ߕ\Q!~s1z­���3#}G����e��
(Ėe�ֹ��Hxvs8�pk#�H��� �%Ol =����Ŗ�'M>�ڦ�>�c.ËQt�'}i�7��O������1R���������-Xa���*`�}��"|?+<%�,c�փ�u��8M�% 
��;_E4t'��8S���$	��=>�h&E�کrc�z��{���䞟���+)���?��0b�����bN-���1p��G\�|d��8�_��S��E 4�o� ���i�b7�e^=��wg�{�'�Y��v% �oD�ۈ�Lr�o�9��A���F���\XӘ��h+%c�����=z��˸b_���܌7��=��YC"֨�:&$��?�¿��n�c��7;�S
Vb��7
,��D(ڋ�#Hq��m��w#��-�M�����t��ī�$��l��J7�5�OH`�Q��iA�յl����N_���5_�"��6�d�u\���7��2
 �#V��ndt��@�;X�d�;�,*G�G��-%�8Xcq�?��n�Cll�.f}7bl�q��z2;W�||��Y�bQ�������GNs����<�`L�F�T4�*����S�d�Ѹ��SX�\��;7�ct�j��/���F�BT8ctE9�������N���������Yü����ߩ?sNa��5�8]�ߥ>�����K�1�s���ftG��3���rΖ�L'K-�<�w\�<IM�j��d`��V7>� �#�8�U��S���lX��XY�N����\v{(�0h����0ߑ[_��F])`�X����+ۘiF�t�����5�6d������w��J/�S��̻���E���H��T�O@��uN\�R���R4�w>Y���4��z�KWЂ�.�~&�0@~�~������+58~}���(�M33}�}�ƭ�D�1�돎�#1NV�NG�B�32�����s�;K�K븟��Ny��-JȞ��弥ȸ����ǥ��U+I����6a	���d���o�ئ���N�u/�+ɼ�d�u(H�_H��Fq��*�T��@	����e0Ā�~���|{h9����G�w������3D�A�� �6��Հ��?�˅k�D�~������]{�S�(��З1n�@��/��f�s�+�-�5����$%,��.ֺm񛆾q�8�EP����{_�@>����2�w��\!`?�K-(� �)"�{:_<{ q-�-�[���1Ϸ�s:���[m��g}5$acm�O30�B���DP7y;�Ϻ��q|�y�U�XG���<1�;ă�"^1�z��j�����8�s���</�O���H����j��T�\�~���ZW�X3N<H�`�/H�$���L��O�?��w�e��A_,N��jd��r���<���4����ˋtq��ȕ��E ��A���H}�Der���s��U|=�J�)=�X�D?��L�ɇ�"^����[oO��.~�f���>)c���j�	�GQx&G�W�0ݙl����數L�£u7RY�a���A��� r��?*Y��C�dVu�ix��'��M�a �~����HK{Q�������k���X���bҥ�XNW�yt�!#P��Q��*6���cs��=ꉡD����G�Iǵ�[ �F�W�~�H���/�K~t�bwO#��L�
��H#Hdj��x����J�sZ�i�M
�Sع��M ����G�@�G�о�@��f^�������1��$��S�{��� ��&%� vS+��1�圕��U���� I�>��jC4T�0z��n�R'��bI&��#
��/7���f���#$7ų-o7;U��}#����~���bl4��R���G�Z�@��m�Hз_vy-�,#�	��P?h��	��C��*���[d�o��#�0e����OE�DV�=Qy�؅��%� �J���8=�c�>=�8|��AW�ۓ5�`��p[�wד� �H�;K�D3�?�����P�c����)Q,��O�1�p�.���T<�Bر��^G��~G,ɢ�b������SVXҾ���?i�g�8��2��75���7��Ǟ���EH\�](%�E�!�q�ϝ�xH����AdȻ�����R0����J0Q�*o���a���R��"�.	�l�ã��c��s��c���a���Ƹ�N�%�h���(�k��|L]5u�.�L5vE-�K��^4���sR;U���E���p^��p:�u��c�j��5ƻ��QI{%�E�}cυ�_NJI��c2@#��m] |�9���6`�ݿ����2�z�ٱ`���V��UU��^�'����ג*f����������
~�U�� &q��Դ���^�	���D%�Ռ݊̕6K(g��ƙ�}Mě���>o$ɽO�x�w���F���i{\�
`}�d��y�g�P�?gi�&��?D"�(��k��]�X�����v�~��O[��2��K�0}�$����lnlBJ}�(f�F�f�C{������=��]ۥ����E��fz�����v�m�ymQ�}�]ߒw��\���8����N>Q��=����w�[VX3�8���ƘE>9�d� �~jiz�R!�\-�iyF�����<Xt�$�o}��<���٬�r9�
X�Q6��z�\��	�63]g�$�N7���O�j�4i�â�(N��ʷ#�]�����Q�8�IHu��$C���"��JT���	~�e�X8��ϼm:�m �V@�iy��76�kQ@;d��
I��S�VhpWA8���Y�u]��3wn Ô��.�X�c�ǷS.���L�,c�E���h��k��(��HP7i�*�&1�SE:ٙ0�|�ⲿ�tW^*0�yM�D�f�b �J���;�+�����4�����qd�Gp�c`�'u�"�i�}#v}O�z�粛��f|V����=�V��>�W62�b|�)~c9��'��J����b5�o������񙉁r��	T�=�{q͹me�r��E� J�b;z"S{5&�q9��j�H�\��i7y�=���G��PB�/<O��CZ�CpW�"} ��3S�+iL�{n[h�Bj�l�鼖��X=>�=F�Ȧv�"$SÈl�5*Hd�xL�*�I�n�{�q�@cj��cޛo	�TW�H�=PI)4����J���tWh�[��}W��=�����|hx�l���Wn�iS3�S�\���#j��YP���03[��C�LC�c�걾�y��Ո��O�+<�[�RN6����e�f9�iҲX�"%�6ɪ���:��A�^#F=�C�;�����m��)�{��E�`����Ȣ��mj5���a���uX�s Qw#|X�z��Y�1�����w��5�_�#��DΦK��6�r�}��疞��z#cd��p�����H2�)]� r���}*=��3?E�dn��Me�� ��'5ԁ���C�@��i�bxI�Ӆ����5�|գ㱴*5� h-, ����q�X~m���دz�������Ί-��a�-��j�m���$����n!	܂��6���6����{����{�o��?����Z�jU�� �37݄. �O�!�r�y��B[���X�[9��)4����,��4����4&i5ġEj��S%6&�Ɍ�U�}���ͭl>|�m�x	�x.E��C|�Cr�5Ou���L=��#�6�v��囷<	)3Vp�iGn��t#��_�ȥ�����K��p�zؗBT_(Sб|��7��'Q�gfi���a�
�f���\�ArQ�� ���+��2b�K[�6'�?��d7 �!�yϨOd#iP�+1"Y�5��<�
�U��d�],*9$��)E~0j����:�|�yL���7�F�5q�������L���������a'���s��^'ֱ�5̬����ԑB���)&G��q]T}x���V�����ຂ�4$�lM4�WY� ���U����Y9��{� K��qE�7� ܞ-�BY۬W���Tg���ha(���@ʾ��55�h���L�D'���v�-o�Y���tn���z	@c��ރ��#�>zT~ǈO��J[@\j~���N/�p�h���(�a����0Q;fG�A���pڭ�b�`̻���`�9�ǽ>���"MYl��t�	D C�^��hA�'� ���t�T�&W2߳NLi^`�W7y��g�?�e"��<�&]L�g��Г�m=��JӜ�9�WP�3��Dc���i���u�im���0�t��7���а���[rF���,��/[����uR*�
��쬺�iTh�,��n�������m!��{��B1;�]������Å]ud|�e��������2�qˏ?�����m���c�M{b��hF��>@��Ӊ$� �"��T��{��Ma棞�wҘ겘���m�I1�5}ڌ��e��L6����Ӳ���Q@��j�F���4`923ѭ���WO3�V�Y������h;��3	�A��?���׸�`�z<�1B��w��9�郫1���7��L�d��26}1?n��RZ������x��_�3�</����\�������W�Q��߾�칗y6�I�@�7��J'�����I��=�F��uU� a��.� g���50֟�g�,(���&��ln���₌��%��v U~R@a�#J��L%w����w�Æ$G�9
vv2\c�W���͇� E�/�����6��[�/���d� �lOA	v�:t!��Q�A��'��xms&�]�4���e1brZ��ە��-����ճ�3Ch���TE}���Z'2��兼|Aޜl�L���a�?��0r�+��ʊ���<\HM7nގ�˅Gc�gc�:�G�V���P�	�� �(ﭻh4̝�3�40ry�4&b`G1Ȩ�j��T��֗�<sޕY_^��{k=���X�!,���@eC����\�g�iuh���"��, ��S���u�Xay���`c�4��	�������;��q�����tx�p�����j	�B.4�\�d}���[�����;��Rp�ɼ�v�X3}/����GP �Ŷk�idݓ�h�	��#��~<�ӑR��n�d��ŗZT����-Rm��pV�b�J��合Q_��#���f��ӌ�T5���*Y���JP��z�34�%C����	��
IKwo��*d�%C�~����3��W~����b:�]���QS�z�"]V_j'�]�luFeE�)Y���Of��$C���۾[%N���#q�4�w�zq��}��r֡ˌ���YkX<v��7��_3�W�9?�8!Q�l�,��XZ	���ν&@e�+�9�}R�T�����"n��p��
�_��ڷd	�K�*����q�aĠ-�j��P���|�sd�C��0Tb�߾XkA;#h������������r��d���0����|�J�괥G�}��of�]��ao�pj�;��%��`�;�3��y�4��M�%bP�부��$G�[3�h4������M{�3��Q�W#Q�KA�w��x��<��׽�
���� Wt]:ro�G��Zl�̞��c����If����=��eN?�b�,��U؄�6t�qߡÎ�q���!V���I��X�#Ş���r�O�WO�]��{)$�?�<v���B�;x��1#O>�����xCm����?�-YA/}��F���vf�;����DG�5�����uZK�o�����w>g�c_�U�~�e�vX��
Ơ�%]�n̔dP'�ie��xNm���U��?ϼ)��}c�G|�B����ݫ�5����#��g$u�����"�s���?yK��>�Y����$����E(~�r=Ww)by��mnq���&Z��K��d�`�ލ:�$�3����u���><�x��JNۏZ��rk����'�I� ӗ��Y�ØG�e>X� �$E>��S���^�;FL�6��5K��\�#����u���x�P��
<�2Pm~�`�p���\����}E�53=��ge�S��֦Xp�*��yg�u��Y�#*�����+�p:�fq1%��k� M*1 6W��1�V٩�v�@L��!A��ӫWd\x${@��ɻ%�^=|T�*�c�<RY=cb��ä���&�����d�F�;��w�-�E���5	{�6v �4�3���Tgl�I����[�f��R������f��P���?#˶;��z�d$d%S���8Mj�)X�#h)����A�z~�}�ġ����w8�˷WYjz��vЗ^��犋8�x0���1$(�S��H0�������5C��)����l��_��Q\��no����|d\���}��X��`���(�P#кM�3��p�t�<\�7|�%�9t��Tu�g�I�E�9�:Iƴ"��@��am�5|��M��%IZ�#`u�<k*����S��I�t離��,�V`,?�HN��Ѭ�Z�A�����^��Vw�L�8;�T���d%afL00���[~�I�j�7EPZդȀ�i}�����;6��9]i�Y��)����hS@�*���?W�J���N�/:n�d/ߔ�Mr��T~�^g|�;t�)�/o���l��ek��(�����ڣAK3��3�K�3����4{��>U�]�r�w��K�1��;�_X"$�Y>�hν7�9����Ħ�!�J�:�!jFE�B�W_��8����l�f:	����5�\��_J$n�;�>qs��.j�7����7�"�1� �7Ԉ&wǗ�*<�s�Ո��Kw�/�)'�i���;U�L2�߸���#�'9$��*Y~����fu��y�`^�Q��G��;`O�-N��Ve}Z�J���a����+�c�����u���%j�1��;�/
N�?Y�+��\jz��k��;~
(N�Cʤ���N�0r�w���H�0��%k-�p�1�M�ڌ��܈}+���a�e-鐹JƏ6�@,¥$����xmEA�É��rs��Y��o.ļßw0v�"��`V����3�p�(5�Y��x�Q*���N!��Z�-ȃ���ԅ�Eq���=��
����}N��H�8>��B�� .w��q[[��o�0"��AE=7)� K1���R3q�S�kN��t0�q��n����Ý�x�f`2 ��Ș�Y���QX��C)��o���s�|�Ѓn��\כIr�P��l4�N�{`�����7�|���xe�)A\E�#$�ԼAE��LN�p��?I,i�:ѴZ(�*��cO|�J����KP%�n���j2���<ɛ|H��ZC^]
��MNfN��%����S�z��L3���Y���rE�ª��cIv��@��5�5��*�.�5�}��J�e��S��LS��d9�ҝ���ӄ|N�&��N�?���Q�|R��9I6��Cp����:�*Z���l��-��8GH��]_u��xJ�i��J�w���;>�� ����.���c�^uc�5�SH���t����3�#�Ss����[����Q[��S��J������G�N2�7&J��lvܵ o���m������GIڶ�Č�΍9�d���+P�6~<0�S=\������(����o��,�Q���$k��B�)4��mIVB�����n�j�����m���l�Ȣ�q�UJN���	埘��W����} Q���ajY2K��,u�CT����P;s��m�Ǥ�p	�! 	�"�S}�"<0���:�4���@�[��S������S��M��~����s���Ȳ����p�J�����6�,��Vil�!��U�|ъ�1�
Dy_������1���� {,��a0�`�)l>1K��#ߩ`�����O�X-ȴ���`E1��X~K�>i:�����̡9"9�UQ��[�ek��PH���4�,��B}�aT8L�N�^#��5tT$f������Y5�w��ޣ-���&b�p6sc��V�^��C��t.F���|�>(ŰZ�'i��X�������X�zL�#&�	��b��̼_�_sG�#�]���@��m�R�W��\�P���W�%���?�K������L�޸��ل_����~0�cݚ��ߩDmDQ��{wP�P��h��	�f��h���� 0�q�
�V�2��� �5�PON���$u��C�o,jin�Z$��ɢ54D�A��B��}��,�r	E��C��H��_��i+2�����g��������{]� [[PA�>X.V+."6�9ڄV�`pY��Hn�*�$I �O.A{[��>=��wxպ�M}h��th��������A1�o�u�@����t��|?��	?���C-m3�~o��Y+|��4��{�lEv�Z�����iA<����;�V]��d�wL��'?g��2:��RC�W$��q%ŷ����F�k:�o��3�8���������jLW��z`j 	Z�u������D���_�.�96���>f�s;�}lU�6�0a�8Cˈ�������"����t��2���?���("�e)_���I��VԮu��/5i%��n?� ��(��$a9Dh��6%����O��{��d��h4�q{;7JROYW�ڻ�ӿh�*�v�4=Ĳ*N������2�$4I���@���7l�y�3Et��?g�`�rc"ډ)�6�*n�$�8�B�W�5�N����0��Җ�W"M�o���1kE��(�XwQ!Ѱ�F}�h��վ�Kk-���kfi�eUr���]��8�Wt�A+�����U�q�~J@����ቸo�u��:�x�MFb�DJ[�@��c�eQ�Z�VS�\ �Z��M7SfL ��*_~�G"�q�8hZ΄����r?O�����T��)x�B��"
S�s���Q�9�7��쳙./ �S���UC��Շ7ض�-w�< ��o\T^)U{�ډ��at��|B����=��%�S�O�I�U8�$��"�}�W6LWT��1|�^;�"oY`X�4�3*,L4e� ��olҎߑ����V(�uް���{!��Xfpq�R�/5�S��*��s>�t����DW���.b�\j�]K���o�͎@azl��z4A���T�2�+i������*B�W���BQ��g�#��w�M��WȪk^dϪ�4M���AގI(���+��_
Z@T��>������i�ҠI5x�=A�푕�����?��zw�|�yV��JTvKh�Lci6S!M[}��k[yl�vTь��V��˷���S�U�U���R?�j#HDf�d �+^��v����@�.��z��"J�D��1��r�11���=_�N�?�����78ŲU��0ކ�ٷIcMV��Yk�j�A�%�Э�~"NrOϯ/Uj�TP���{�]�����\x���pv[/�y�a�6s3hI��.��.�����N[C�# �el�=��j�F)�x�d���
���2��@^��J��w�5%xXz�5{E,������'V���M�|hK�L�o�ڑ|[�M����׿���'�&�\��qz� ��y2r;7�mv���ə��S>�?u�7�[�tR%��js�:�7��w���׉EЗ�܄eH����&�{��U�j�}V|D=d7�`lkVM���M�����:����AH:Oz�R��k���ү��l�jgG3Q�	!�*����}��%+"���F�݄���U�=��qN���1�{�p8�y��c#��{.�u�}.3-:�-�'��_+w�]��)�=�{R썍���2�=��?9"����x����.�<! �o���G���jy���s����a��L�<��0�X7=��@����A_(Ǎ��P�����n�7[�A���f�,�"�͔�"�d%W8�T8x���ڶ��뾯�^r���ϬxJG�	J����P�o�	�՝��˖&�#�9e����7���D��[����1���jl��˪��2���I��>x㲦���ꯨQ�'�:q=Nr���$��̋�hog��\�Qܜ�I���VZY��xo2�i=������L�	��nȗ�� V���C�ߡɒl�+Щ՞��5x$	2�ϙ�^�/I�D�c8����7B����?0�����M���!qu�eנU�r7��򱽻Ǝ[��aA�cF��hQ9mQ������5f��\�J��w��Nk=��E�OA)
uy�ls��s����v�u�]l_]5�J�9_Q�r9�PJz�$�G�#_�߯u�ܯ�uv��i�s�8����8�]���ʪtݬ68ޭ!��<�I�������[5����	c����}~~��kV�S�����A	����aݩ �xl�F�����3��D�[H'�l6�y7��V�w �((/b/�9�����D�;��(��bSh6�d�OL��T�U��"''45�l���!(�j�gf��4��\������xbWX�U%+���۝p���7p�@u�1fRk?v��@q�|"�!*���jʗ`�������K���R_9(���;A��X��m2�3ļB1�n3}g�xAZ�z�i�S�!����p?�:��Ջ8n�.h$���%(b7�Yx!1�8S�N���gz���!i���`�?���~ _�/��5Xb}��l#m��AJ����R�L�>��iS���M,.q|aޱ�jk&y&AU�x�s�%� �E4;=� 3���ޟ�uZ���D�dKva��х�H�h�=cn%�%Y$	�!�t�I�\��W�CE�[	n6v�n�����5���U��Z�NĝI��� d�~���W��]-?^�<r���s㝱 e^w�r.[�����-n@�C��ę:ru�"��^w�]���%-E(![Lu����HS��9Ɗ��e��U|O�U��,����_)�5���JgY�GU~E�ݩ��`��-�{�����<j�P�k�#���ٿ��O0�(%����3�v�=�	ε�{��BMW�/F\�c�e
"�&A���,9�G���ȼ�ֿiE��Ya1�06�Y���?	�3��r�S�G�?�O�5$é*Z�:���M#Uls���%�Η��ܟ�T��(,�(?D�ƌ���Sh�0�[���������__9�~� ?�j�+w~D�(4T�g���r�;b��������K�9�+����p�?>��y
aV��
��q3��L��z�F����g�t��ӽS�l3���X���b���.;\���[#0���sV��=T'R�-��I����M��{��!�j~�XVyl�������
�0K����u.FǶ�}������Z����d��%��eђ�zvڙ�Y�Ɓ9�t�d�8��S��۷E���w&�>t\l��yf,y��1U���uwڹAJ�E�Q�UM��;�݆	aB��NE]�νa����	�B�� e/�A�ߨ�J���<���=�0�2U�29`�^�9s��pMu<�U쾻D[���ժ�&)�z�|�P���N�w�s�� ��5��H�.���g7�oc������,������v>ܸ�P��F��ඕ������h�u/�t��jm��3+�9\��?��T�g	@�yX���q=j��ޭfd{/,���B�χsz4 .z��2Y�keo ��1ҋ�'1`L�83�dɜ�D̠��]z�i��C�ˋH��>C� 4������S�[�a����ɸ�iF�����.`'h=AVC%���B`J,��W!�@�W�@`�d��������K@m0HB�*?���2��/-ӫ3C�B��FU���S���F+��&$<-Y�S3��pbf�v��	b�}����m�a�����,����j��>�.����v�yg��Q	R����sڋ��\����G�BX+e(c��K�sM�+M��c9ABj��>c�'K�͔�n%����S�a�.Ͱ�G�A�N��פB�i���Qу�ta��J���>�ͼ�����6��`\V�\gɯO���9��aP�řC;�FČ����"[���C�`RJ1���{� {���[��m��/ow���@gKvCzC(�Oi���_�� ��|$����D�h	���8�5�1��T8,�w���q
=�Uƙr��.�w�P��Uf!"�j#�������i�/�����)��0R~ ����'+��:�S���3}�*��-�a����SC��z��2�+�D�&�{l�'�0���L"7�.9�a�M�33}�V�42l��]�6MA_����hˤ���0(����h�<�/���T������ރ����v�Aʄ[�΀=��&�����Dc�{Ƙ�@�]ƕ����G7F���������yh�YA�FF~A����ek~3k� ��)~���~���{�O^�
��2dZױ�*��d*����&�T����c|]4�*L�=��J9+�ds>��)�$��.HH������EM����T�拆3��hY�rs�B�
�l�����tO �>b�����F��l~��u/�������}W���;^���[��i�p�\u��B4�"Sʖ����-��J�{1r3�,{Ǝ��X6��L�ݎ�Q�8�?�r���zz�`���r�7r^@����>H�c����~LH��G���{L��ʬ��vBVD�m�|��
��P��Xf�h8���G�� �5� �.�Ed��]���x8}�-%�j�'��qޑ������ެ{��%���-Oh��n�Mǭ'Lr���QQ.���%u�1�	�V��aWtO���`_���^�׾R2�C�%@�j`�u�cf��άs�n�Bg粈K�Lm��5����q�eR��%BB�<#s��#��)W��⨘�$��d^&l`D�H,sa����YL���\�i�3�[��ӥ,�VU&��V'JM��H��bl�Wg��HX�����S����1]�M�Sz��i�8z�A ��X�\|����	v�4�h'O=��&��>]7�%c��v��V�Us�W��g������P�}�ua��W�P(�:(�g�<�����:f:�V�����f�6���ILD�ܽҫelI���
�ى��?����ģ~f��H��-. ���A����g}�In��U�<]VH�@Y�/�p6"��^��r��5�H5��ռ^[V���/��r��v�|��7�qv�����X����p5c��mA>*�7JF��)��L�nXY�LO^M��ߓ��ד���h����?�a����ה�r��-�8�B�h4�����N!���(��%�D��t�%g���w��Pŝ�5p@�=���Ԋ��7������E�\���}C��⅐�a���@�K_z�K����DZǏ}�����_�~6p��4%�s0P�S/ �T���|cbEĦ�^Pm�����2���F�]���P٠-��X-����=ƾ}"����J`��{*6��h>���Zd��������e�r�pv�I�4����3b�X)���
����j���x����xMl�?fcK#`��*k�	�®;���h�A��l:��~����jl�
.�0��c$���ʱ; �q�|t9�G��
QAT�M���n��N�˚���o��Ei��}�,�n�Lr�*gEMm�S�F_���qA���t��	��֬���:7w�`X-��"՘�Ƨ�����(!Wx"x��v}�����Z�.�/]nƯ������_[F���c�$��a������'�4�P�h~j�V����i^X��&��.�5�'�E��U�/��h�o��N����@��Hm���9r������6ժ�R���Ӕ(4����t����b�J�8f����#o{}��1��'��N�0�����;P�lw��]�&��{���7:͙�QG3ʳ�h1��ҁ۱}�ض9���E�b!fO��d�4x��������W�g4���Ġ1ߧ�"U,"�r��~}h�i݋�x,?�'p1���"�scF;�-Tz�
ߪad�n�˒e ;�Ef�m��^X�>̠ܸ
��%l����`rw�M,���hkf��yT���w���U��͜mߜV��e�D�O.�C��J:{��Q�����<�`��D�����S
R�3z_��Q
���J9\t�����v�� ,�g�����^,�{Gʰ��!���f���h��M���|Ψ��䙢�^�R��Lv�lnQji�m|��$[U�	����� ��j��ޔy՞^41����:'�8��Ц��n��[�1_g��R��r*�,>�����_��\�<s<����p؂3!x��7��#4����G����Ҁ�G{ԇ09��p�C���թ�}���x]�޸���s�H�;��ư��6�8�^T����[���-����NN�˜�X�z�NH�O�X`e�1��*ק��N���_$�&�QCէ��}��t9\�YO2S7}7��8�~��J0��x���u�8<�Ё�a���Hv@�a���W������G���^�r���8*ƚl���ࡦ�Y�}�?�� ���Q��2�[/X��M����%��+���z�Ji�+@Q�'������3S��?�duĘ"��t��W�iJ��m�ţk(-Dg7�Z7�.enpL����,2��5�B���B3�A�P3�ȸ!�6-��b]�S'��rU�>*?q�<�T�\��y	����y��*�#��������?��eJC��;�3Y��3�6N����5C�*2�G P���T�g�@�w5����$��'�bTX�a0�Z�R�*��\F<m�\��ڛ�)j@���
n�ʲەO��b�ҹ�Qg�Zü�@�K�\�} �8y�� `Q������bB�� �0qgMG��V���}'m�%'�����+���ۣ���`{�- @N��
f�y�W`h�)��j�<�+��,a02P��\�nAn)JKL&�]����D���ІnCB c�x4xL'����M��}
�M��\0�J�7Q���rC��ór�H{.��<� ������9�0N�	`�B�����O]ȑie������8_��d�`K��|o���Z�!ǘ�� ��N��rv����[�ߴ���/{�t�"�X@R KU�&�n\�P��9.N���,�&͌7t<�k���L�4`�:ہ@�|�*Wz�'i^���-L|5��&��卌T錚9�3�n�(���__��N�&�ԝ��V���-'���g�K��%̞r�L���f�Tm~/�d�JǬ�ǨKRc��E�a���(5�j���$[1ƨ�֒ua���B����1\���Ćʎ�O��o}��=��51�6]r[�u ����]U�lZץ-�86$���K�L1nK4�����O*��ϛD����3�V��7�9��y�92i�͆`1&�����w/t+�9 �(� :�~�z�q1X������na!G߆7ɗH�$ I�T�hr.Z&�=���D��켰 LG��i�E��i�E�dq���}ً��m��,��b�^߇��H-����'Rs�,�ځ-��X~�g����M���].�Q�&0U�%�{3(��5��RLDU�}���|_�ЮQ��ab���5���x�=�ڕ����[+sIrb����͈͕a8d�A�4�!���7)������ 1Bv�y����#_{i�

�4>�cGe�p6糶�5������
��p�\�R�+'֏��~]z8���"�����@�m���uk0kX����\~Q�r��Ѻi�_�lS��FF�Ǐv	pЈK�sa�xB�[�e-�yA�N���Oa���L�n�J�τndMoJQ�����O�6Z�J]���?M����d��%*�B`J����'�	g����ml�L\g���̙y4B^&3����'b�9��h֠Wd�P������;>���|[-t2RVE2�na^�R4f�"���Q  nG�As���n@ÆB
���%��Q�;ߙ@��zTU�ή:a��uL����>U*�yf��fŖ);5"pM����n%M
%���e7���M�wI���W:�twD�g_��Ժ.9[_�b�_�e/p�S��5ߝp�,��}�>�_P�p٫`߾y�'!��VB��h���)�;�GޓH"��~FUU�D����'��K��.@�>?21���s�f ���� ��๩Fe=���6���<���Q��FȐ+:4:3�ru����CńH�����9#�^���ey�PGB~� ��Cq�G�W+���HmE��v�lf�q�Q�������V�xNɻ4��&�S�L����cs��~{�.p;G�`�׸��['�Y�9��IBZ*Il\�O\��p�i4/��c�5������
ގ��u)a+U�v�_���ի^t��C��9Z�e*�[��;�����=�kIωP��H�V[Y8���%Ձ��]��$ ���?����(��ʶ�\,ܰ�j\�,54U)4���ά��H!�Kzs˧p�о����������c!��`�q�	� pu�o��,iB��VA"j�1�~�9�08�@X�}$wXZ�����`8I���.Ă�|s������  �uj�PE�֕ ��R�������1|�� �!�9����;�-o����/�6���.S���Ru�1��=7�R�A�Ŋ]f�_
�Q(M�o�C	��i����� '��{����(nf;.錰���<��*-t�;G��C�{�=ƌH%�k���'G�"H<3��A�;����?��X�w��b"�XK�c.�8�ǅ��}4�vw�����S͒Pp��K'�&�O�sX��,.�(�#�2y�EP�DR5l��->-U��Ozۛ�R[��T���|���jn;%�s)-�[�4�"����
=BM$6����`�g�(�*��7�NC�ZA&���\T6�]�ϮC�Z�hG�r6K5�<RIܚ���z��IJSU��`+��٭����? ��A�^����|ˬ�y]?��X��Ő�+.�D�!:6����R�,ks��)�C�����hq��!����6 Ma�h�B7���z� 	�����C�?�ۯrڜR��qߨ� �FC}L$4�;�|�w��~���s��:������6)��1Z^P r�Ĥr|[k|[[����3�#��'�q��a��� �;��`:��H�vg
{p�ly}���K�Qxdx���а����HI�
�3��K�-E�Zlzy���۲/�fD$��p�/U�8�%Z�q.�J������6�s���v����G�<�I���30p�\�i����!LEa�Ԇ���큦k�����S���yNO��R{�����~��� -��w(���t	��I�睘Aw�ݛe����t1���:Bj�u'�ƣT[���~f-��� ��{#>]j�s8��ߍtV
����V#v����z��;�� ���MQ���2�I�����
�aPf��k�S�ƛ�&�?�;�:ɭ��i*(H����@�J����L�ԾǷ��yMx=sy��F+�IA��Z��;���IlZ�z�wU[2I�Fn@ ���7e�܋r����ޏ�J��6r���Gz���J[*K�,�+P1}ڌ]�������S9!7��aOh���`w�w�|�7C��}r��ԴA�����IJ���Ʊ&
yJ��2�ZY8�h�%�4E�;02��1w]q�`�KG�'4��	��ʥ�0�.��o��Li���9	�@����:y�a��FEaNk�&aJ�]��m�o�����$�R�$ 1�����t��k�a�q�&As�}�����T����1�7��=�� ��tWQ_d�b��{5��O��k��'9��|�A�F�}��>|!��ݟ�e���&�h��:����|q˪231��1m�9�=��ְ,n�Я�h"^k�Vv11��@�w�Ǝx��D�5����-Dsr�Vo	�W|\��r��b!����Z�NX���Qf��Oj�4��aeWG2�ע�ɋ9�ߤ2�e�����u��J��~U��#�"�X��׎����\�_z��_V���"�J�'$l�Vh-t����w��[ʾMD�4��y�� w�9r�>p���`s��?1��a�k����eQ�ɟ���L�^��ރ��4�3+7_�!�%>/A��8a�1��C?�h�kr�ȩ�6��;<�6�ޞ��y�I�kl[K�_�6K�-K/T{��ʋ�DЖM
׆�wt_��ű{���&dl���t�a�?8c����M�p���#�=C7��K�o�pv$c≐K�T�59:B~'D������ ��Җ�]t���Qd���\=2'P������(<��te@�)�I��ž��J�Lq��y�.�$������5�#�NXv���f����:o�׵�Xܠ2�T~Б���������G���4�fY��X9-�va�
%ӆ��3�"
��&��W���������<*�d:�j�'�&�WHp~Ac!�i���:42�vH@��r��)�����y���C(f]b��*VO��ψi�ؙ$�B_���o�E���ɞD�'{(���φ��o^Вb�T�K#~壟+�ࠑ�8��=��xp��z9^��)H��(9�Q���Xc탈,�A����Jn��ȯ��!�5�@h���
�H4:S:U ��8�Gj�4IA�v#ϒ��{h!=|?�(�HH��g X��j��V���^;2�Jd{�P7-3����^�O-:�o��ۖ�)���8;���.r�?b�U� ����"�f� �b���fF#�J���eWk@Ĵ���L�M2�(E���8�K�,,���ߠ"Q�˖crai�T��*�Å�B[�	^�`�l��)��/�r�@�`���9en�8���b���,r�����C�H��9UlK��a��$�U��^�G�7������dK��v��q�r醡�'k���=o�y��˛�h��!��b���t�-�Y� ��*���$�--,$�S�� �1~D�7��;�N)X�zN��X����vix�JG-��êݧDKU��<	Z�������@���� ��*H�M][���E�yq�nf�^����QJ��t�#&2����?������o�5��C/4���%4�L���~D|�l����5J�C>��E��E��5�����"�P!�:2��z��KiiH���Уu�儸|d>��s1�h=FbòϹ1��$�cu���6�A�N�����!�ֶ4Q?JcM44�����E����xFBX����>QZَ&%�<v_E���%V2Z�^���ѝ�9_p��>�ޣ���ՠ��8KA]V4������Q/b��f�7bt�~��2���6���| �`t�����]?��"E������ $,���I����E6I�~��l듚�sX��o�B�)Mͮ���r҃"�n��L\�'
���)��mh�8{�uҚ�y&]^�����_M�f�.�C&���'BknE�ؑ$E��j��? ��L��#�jd-ރ1r4GE>�����,��N�j/%K��R;��b��>sK�k&��_�w����iN�B�.k(P|�ULS�K��񛷗���;�ϯ
jh���!�+�@�=��X���h8�C�e	$	� ��r�b��5�I��l&&ւ�*��`�o�x_C�R�k��\�7����	!A��ɷu�[�DE|H<nzl( �!��9��Ti�;r��g7�'����d��_�^�<S����1�Ѥ=<b;��U)�6�F�M�d3��h���^�q,�b)W��=�fip���r�"b���o+Z��6?H|_Q秔'v�S�^�	O����������ھ �C�t3���0��t�t�P#��1�H+ �)��������>�Η�ᬵ��]���:o5���U_�)�hQ�[PJz�Kl�al��L�I�F�	�q�]l~����0���E�zF�}�����!ߨ�\'��I<0��f���S~����p;6"V�(�\�r��_]���;J�.RÆ�{Z�/��r�������D���+ƍl�c�/��������?���ϰ��}�K�CG���*S���0(0m������e��=�͗��_>)^�E�V3��"��rV����z���Or�J�5�떺��Mz�������䮂ZS�
s��:2]��\�{%��b��K1F�J0�Q<F֤;���6����ߺ��+`�z`l}m3Z����Z	�gɡ�V���X'MR���h-��\�&͑���+�x͙���;�G6�D��XC�\"��KV��zDQ%2���e��"ۢ���!)�Ql[�AZ��'z�K0��Dh�|����\	OZ�n�l^KU�:�m�P�C�Ѓ�Θ �|bf�CƓ�C������U��C)����3M$ƻM�L�7�d�8�g��(b����ƃ/%�C����қ>=� ~���ϒD��>�]; Q��.z�㮾������o�4ɌiK���}�UMq�S����p�{�l�%y-C�]U1�z�V9��ށ	aW1}�Vbd�+O�����+�c���,��V2��5�0�����'L��6`6�Y\ī��@bB�=��W*���C4�k�c	,+}���{6M��f��<=g�+]�]骉��tݳ��[$$�]{�s/tq����kȴ�[i��iF�Y���s�_��x`����w���=n��NW k��F��dio�hz
�Q�[����U�cj�w����2fe�ph�,V�H������X����oP+
�(�PĞZs$�G��r�LC��̏q�c_U/��*�9����6�O��[�D�
��4��'��h(�����h�b�apQշS�g|�D}-+�lz��M�2rI��5Z�_�@d��i�A[�
��d_o*L�3)��Yb"�z��&�x�+n���zԐ�'��'Q�ǊI�K�2]f|�S*w��t�:������9���ߓ�%�����zjb��IcL��\��̙Ad|r��Q�.�M�۵i�W�B��/(��X��H*˭o����N��!�7�8Z�P��#��U��A� q7��A���b�M�#s1�{�	�^`������5f�Uy�ׇ�o��-�pX#
V��ўR�F��į>kD�24a^�{���F�c����X�����E�ײ��m�vm�>�M�f����#�+��dʡW�v��5,t�z6Z^$�����r�3�\����pUy@_�0 ��NC�u�(��`&��2E@J%���(/ȋ�.�t&�L���}�03�z��/f�X�-(I&����g���@q�Ԇ��@ާ��������t�1���� i4���ݶU�W��3.��#'�w8~�^��T�f�e�2L���!���;�mqU�RW�����>Ѵhk�x��v������:�&�P�5�Rz�v���0�A5�m	��JM��d)�K��H�-�!	'����z,D<�DIޮ�׿��ݐ�~���kYzo���1�-1�u���gJ��E��c���*��,S0�C��եi�L�4B�|N"�֔����c�{.����~\Md�^���0g����U$��4�0UG�"h�H�z,��֦�D�'�#".��?x�5_�5��"Jo�n�h25����Z֐�p�HB:]-�S�ͫ�4�T㾍�LjB�����u�Ҕ ��U�GB��К��
"������6iɄɻ�s�k��g;��f �A��z��;�O��"��3P��l���UN~��*�N�#��/�L^�ޠ��O#�K罦q���헿�PG�GKkY�?bk�jIhɏ��JDoi�!��h��s�GS���M)2�X�E6��6	��ucP���6M��� ͣX��%@��D}H�B� �Cf��s��$�Qi~����@�#��4�!T�3#�}Ȏ':�~�;"�vѧ�O.
^3�'�H��i��+%h~���q,���A�ˇD��6\�e'7�~����c%?�o�	�1{>]��|6Q1��A�D���hAD7��IyS�BH)�zT�,�f�0��a��w���cû��M�8���}.�Ƴ�y��0'edp�K�����y|�7#�;�������l��U 2M^�YI�;\�^���'��ٛLj3l�l*1�j�����6���y�Χ�s*d�]B��곁/HT�v�����)w�����^���:���Q�����������aFf[����C1�=�N�_���J�M�ꕔ�����5���e�YPH&���_q�{7�,2�����"���&�����3)T�Y�ꝅ�y�(�����w��ҁ��$�����T��*���p�'�U��*���$ +�8�ϡ�Sg��6(��	o�&"�B�&��@�m=�����'�O族�(�6x�J�;��Q��etu�wa���Aѷ�T�ϳ9mk���l���o�3���-�#x������<wY��à��:T|�p<��a�n��o���5�uG��,^�ڮKml�O��$O���0(\���?�\xT�)�PIE�w�O�ǐҹ㤵|����\�3F�;��� �`ƿ��@7ֻ����(�|��j�Z=tRT���趭s9!$Y�H����u��`�V��b���	���H�g[*����e�����ƨم߇w�^��o7d:��Nd)�u���nS]�[�a.�2�����Z��V���a�e?���io�r����>Ix�K�54�cY�G��˔<�??�#S�#=аpQ�V��/j2^���c��>�7����˿�.�xZ��6�]:��~Z��W��������H�����N ��� ib��Ve�'��Du�$6C�zO��L�~�#����������g$��wSM^rh�����O�&���l>i��tH�[7��Y�Ue3�e۸a�F(���x��OR�[$�k�s�1vogxv`vt����3SN\������}I�_�M�<�%��#���F�r0���b- ��|ñ�=�,,��FG2��m�H�N�c�ۂG��u��T��U3%̅}�#��"A��q{��p�檕��|�7.Z֡~fx�s�rpCi��z��!��a��P�f�"*��A���s���]��U��"$>�I��ߒ������Mm��/�w����1N��x�(����{�*W�巯�Z-���
t8�]��Ԕ���tY�����������N ]��6O�% �Ρ����(�i�*2�����Jb�/�UV�ߔ�1E)o~�����\��z��o��x2��G�Zz�}�����[���=���A�L�d~z���^n�<8yDşz؀ݷ�F�%~�]�X#��S�@Y�|Է�:�q������(?"�Y��++���i(},�an�D�AD��Edԏ�+B0��#r��L �	��C�؋����ɿ�Cp�[YҮE-���ǀ���,�JߙL$ h�I����ͭth�������j��{�G�?�MdF��Q/���j��{l��S��NS1���2:�x�bё4�:m�罻���P��@��˹�#��RB�pr@b�C�F�����$�s�ϊ��N_G�8����v�Q�ڦ�1ˏ�^��/Gͬ�g�q�=e���4�hx��m�6@j�s�g�-y���jo�P���� �f�Z�m�D��::�oZ�x�[(|dQ���Cب�n[��G��q8R����G�7C+r����&��-������0���fw�"$6��T�o73��K~'!�h k���Ҟ�1�������M��a���?GM�+���$m��������pa���/r{�p�~���~tQ���z�l�oKN-�����Lj$��2"iV*m�kL�mo����(Y�"Bάu���"���}�2�|6�e�P�Y�.�pX=CA�J�0B�M����͖�a1������ֆ"�#G$�F1W�O��	=^��5�&���������E4Ɯ�d�3��ګ�}
N��o������|�.�l�C�%������ѕ���-�nFԅ>�����}~|E.�PU6�:�p@�FWO�+t��*~�,Y�X�צ��F>߰oY���E#Z��Qd�F�ʣVaJ�����xL%^ ��O8��������C�Z�$V���^��{��jZ��M�D���~����8K�&y@�E�c���u�<���y�Q,��rv�ǮFb`�ɰ����p� 54�PT�l&k@;R�)�Ee����\9Lu���8��E�/�K��������$"#+�6��U�͵8��-1>u�U�ҷf� ���f�b)�s 5�]c;�F�a+�Z*[���i�G�&%�z�{��e�b`<Tj
�F�ō��z�$3�h~��L�<oq'|Z7�����~��k\���-*?8��\�V<_$��k,�`��,?!��.��HS�"V���m�ŪJn������&C�����;�Q.�PG���	u�ޚ���:�c�b��<�~����3��$yj���m\������|F!�'X[�B�I�Y�C��������W�&���ȱ�%]cQ)%R��B�J��k�wT*M1_Y�,.FUS��H���p�o���|3 �3�ep���t ��gW�K���*�|,���^g�������;n"�uX�������*D�ݛf�g5�g:��
��4b"E��Y�\�3l�%t��cJT�rf�%Ւ�K����)O��O�ԉ�˲���U�̅� ��9����P�-�ɟ��j�q%$��~�2��Ë<Tb.�u���u��-�l�!;�^��o�)�����{z��r��_Q�0�w�Ʋ�ʔ�(J�L4�>?�����Fr�Xl��SA6�P����[Q�1��2����Qw�6�틎���=�񲬛"e�&i��R���lk�c?f����*���_`��q��it�r��Ŏ����۲�I�&,�����d}���]�"r�{�����1�1l��B=���I�F�b��B3�0�像F�����X��Y��!��<����o��b�V�ǀ�\�J��}���\�`i����8���3V�#9MEK�d�5��	=��k7�����;�F�x����<�|Y���_���M�%�e����:-`�W�\���?ǃ������w4tР���?�_~Ka�����K�t�����U\��bc|&he�֢?D@'���Ǥ	�� �V4\��*� �b�XK�i��_)�DʒtM]A�ögk�%�Ĺ�P�*;�l����.�ς�`�Z�Ev�K��eT7�hj�Y$|�P���˃�hN�vU�Y�]�>hp��qM���n����SypS�F��������c�zE��I>%T%�B���z<�����K����D�Q��o�dO�G���jqЎN��f��(#�Dse.��B��Q���o��]�٠1��T���h��f��_�U������*�b�o�m8��k}z$pŏ@7���Yl���؊���٭�L
��~�O��U9i�����e�U%Vяje��}�ώT�iHEX%ڻ=�t�m���5 ����IpT0�;5�)��e�h�Xk��N��iS�����Q�}SF%�_��I<����]����du���e+��s����[`�*�#&��цԩ���j~��W��������x��44ܛ��qW�L݊���ͫ�S�|)�Qd����O���������?jh�Ah��W�����Թ�OQ{x�����5rz��|@ �s"�.>��T���)��p��H�U�:S�"����"�\̮�H7���Q�\�,�j��I����p)G	�0(����$:Z'toq��-��5+(
ۊ"�b
�4��*�c�QSiņ͛nݓ�^
��J>��+�1�:��������-�x�X ʷ���s�~��ͩ�gqp����+�y4Ɣ`�4�%�(A�,��ktt�LcV��|�j�#�rx�T0��}I
�[��T�PZ�I榌a��ū�ۓ�j��E� !������'.OB@��J�a�T4��mq�DY�ʳ�SG��\�^w}����P*��|�G,�������=��#W��_�J� �͏�_x+����%��ZmYx����V��EY��?�n�	&�:!ws��y~w���>UK��<|9iᏹ����z�k:���W�w���:)]��Ss�q���nm84��mI�$e�[�S�d��4񢁬x�zҷdcQ���"�?��a�sb��%���#M�?�e��K ���8���*
����|��'�P�\V:�_�Y����)B�U��#��D���؇8*"?I�`:p�{�����@�P�M��8BM"n89g�R�g�*s`�ܯ2��r�l���x���/��D:^�J<}��	əB|68^N�W�5�ܨ\&q{0u� 2�������G�H�OkkEow��EX��L��]�ӓ����f����ί#�.�p��3ˌFH�!�<еG�d� �3�܈1��}���Vd���l밒������t�Պ`�7%#�S-�r�t�'kR#�AX�x!���
<�W����:����t��ړ�q���`�6k�Q��kt+�g��<x�ѕ�w���,�<��f���c?��jK�S_��rƊ���ã�MV8@=�����S��`C8������	u@��i�9˿ v������H�h�~���w�,^�Y�)�i;'�xQ��	��|��5v��ow���l��]�ki�83��
�oh�*�.^s^j)]�};�gw��MG���0'�������~'b%�>0����=�a�@\�c���]�ٖ<���U�w�[�b�`e�뎳�{���GeA�����9	���b#������⢽˫]EH�].:4AD�w�#Ec�;&�A��o�� �񉬊	^�o`ַm�7�4�?�S'/Q�r��~I��bH�-
�(� B���"���{(�ج1�_��Zi�z1���*����/$��Y�nv�D�=4�W�+Cߵ��A��߹��%=��Ϻ(Zx.2+ Ə��xH"o�GP=�� � ���=�7K��ZHy��p�o+Q{n����Bcl�f24,���3_���+�}����e5��/�3Fe�Fmk����8E�����
����p-�Q�>�������]6kIά�-�}�|�U�ֆM�S�R���~��
i
�?/��mK_ݩ."�+�Nx���r���2�`'F͇®���g�$���&*D�/��\�i��7��)�h-<oWf���(8�?�S�"���M�5mN}Gt��^SL��� �#��
�U�?�t����(�X��A�Z�@�ZQ�4�y�zp,���87�^�6��:׽�F�1���[�T����gD_Ii��Ʉ7QL�����v
�-����_��;i�����<��ꫮ&��Ʋ�;+�w !�Bt����������-w-1f;gzGX��A�o�ʞ3
��~�����[ ��˅�4R���Uz�Q
v(FI���;!0G����z��ϔ�@���L;�����K{�أP����?�v4�p���P�����j#��)m��/5�H�{K+����tk'�[�Z���B�|E�*��ٶ�K
&��Sƾ��m���JVAww� �O��ͷ�am.�y?�S�ɓ��@���Ƙw� ��i�F+|ٿ����[Tސ��J�{�~ؖg��KV��&O�L��ԋLy#dߊZ]�p_�Y�����d���~D�6���%~\���)
�����'����\�-%|1�N��V�1C�ht񋢼��d�?�|#b�I}��Kߖ hO�P�c`\.� Z��Q=Z��Np�j��T�/��>L����!�ȓ��`ҝ�=���u{F��`���'�>v�A��L��:��lPa�O�z�To-l˦I�W{��($�[˧w"J�Odj$wx��L�=��Aꢁ� Oa�(Eg��C�]s�*�&f�wh�H�����:Oy#�Rp庉���5��e��</	a�I�]<�p��_��5��\����}�n���v��ր����1��~����p�k����a�3�6�����g���	�H;���V�����YPWD47��R�MN�J�mD)��?�7���@X82�C�pCp�������e%ؕA��+���cs��X�c�㤈фȴ�)�RC��*\�sk^S��∛U��X��@)_=��o��_'w�=F�,�+;��Mtt퍱y��uI�R��j����USy��:{��^e����
:���q�r_Y�r�T��Ɔ�KѾ"/��r����-��ͽu��Y��|��$����N��)ӅͲcl�1B�TwV ѳ�,�Odr���X(��}N�7��<1�7ӡM���K1�,[��;G�v�����9KO����D�M{u2��몌y���ɟ"�y�ג�87������GϨ,1�bE���7ź���_��5�~c�ޮ=A�����d�m(�kѪ)� �T��!	Ƶԑ}{���!��^�F��R��0x���wV�����x_��(pƪ%a$R̨�Z�fy�u�k3n�dx�64r���� �C��O�F]|M͍����F�a���ԛ�q$��if��J>�WJ r��2S�a�j��L:���,O-fυ����:���잓u��M٬m��:׶O������^��4�5:4�J�o�C�o�$o�HW�Zi�hvq��t�V��-�?�ǻ���s%�H�R%�.`�YbT��4 �p51,%�芒�L�H��%B&�B������5zvw�=�@o\��I��*�A�r��� �T�b�QҲ�#�̷Vg���`ݿ��l6�؛V^R�~��eAf����	��wm��p����&&A��<Bِ�hAQ��v�����>���3��:��4�Α����U8���ϖP�|s�'�aEI ������8�=�Tu�.Cmj����`�ԤcyQ^���G��'���e,��I<0�#�!u6;i�Z�,|�\I�eJP4~�낑�]��q�f�.��d&\W�7G�����q]���q!���{" D8��]��/וA���p�hx��&Ǿ�s N ۲~����w��,�h���)X��/�x)�!|��l5Ƈ @�83*���&_��@�Fv�(��<n#𖎸�Nǘ[~����p�@��������R8�%ݖ/F��#G�Ғ�I֏2c4�(XѠ�~�aI�M����d͐N-�ME}_	��<����a7Z��6+��Uh���1?f_�	S���jR`ex�	`���-���Ln��k D��/M+�Q(�o�N�����HF{s�&������+m�F#��I�0h ���R�hR��{o��_d��7Q�L �$�4m�0��ݏ\�� �/�R�s�c�K�%�Բ&8p�=.ϛh?�\̯`٢!'{����h�s����؞�5�ʂnS<�h 7z�o����S����|��P�q��!)�C����_8!n���z%��~�X��,A_����,m�E��UZ��H��@O���n�Uw�!�S���s%�uG�P�9��&g쨚PX�ގ�g�m��l�X�F�	M���:M%�~�U�s�R���>�mس�G������5⮱�07m�/pr$��f9P��FQ��]�D�?B-!��(���<zG�ɱR����k&\��J�����H�R`'�-<جz��FU;�_�2��ah�`x9�L�*7������DC˛����jv������'҃P�yH�ɺ�n ~r�Р	��G�AN��q����Knv�]Q����j>7��@�'i�o�I<����zI�O��� �9���%7#����񓜂Q�ک��D�.�zG�=�^�[��������xip���D��ߗ�35�x5��x����R ��������nu��g0�4��`�P����K.m0����A��^l�c��B7Y}A���r{X��T�WD{z���4؋#��g����LC�S��-VA��j��P�s���� ��[,-�<쨬؁����z-n�A�����\�3cqm�o�AS�#��l��,��OBX������Ia����mO0If1,�
�!��"^��7�n����������j�"�]he�2��b��e�9����|ۯZ!ܧ��n=�
��G3����%�"-a�&��ޒ~t�~&�E~
�������e�M匡#�N̻7�����q�X,�=�D ��R��ìcǁ�Y��������kAN�zFcĦ��:���k���0��ћt�E^y��i��M�Eu�������8k�p
�k��TJ��Ф@hB�?ÿB�����w���^��\���27���dX�3̩���<t�+�+mF2�a��7\Ĩv��Q����'�kH�݌�Ŏu�慧�U�EAZs��^�P���y�����N���P����y��@�2y��.ɀ�8_M��f&�P����셤��b�G��3���/��ks�U�}��{v?!��Q�FS�%e��وåJ������FR��Ѱ7_�����~8�^�D��DW1�<`�r�g�y�}���J������=_�FOY��l�˜6����9�- �x9A{�x�_Ӓ*O�خ�����.]Х
�[�*��:�KMјw�K�,��y2�9���X�l�e�ES| �J+���r�ä�v�&"^��O�t5u.D�DZ�JI���|-����2��W��OX�e�<�e�!	������Xg�^ &L�7������*��p�1E�
���6�\�v����D�1��.�3�UW-�B��EQ��䨴ͥ�/�+���!���%Z����q�	8��7��NH����W�؍D C����^���
�_D�,Љ+J��6>��`-��F�ˬJ�6ev!�1^�����K�w	q�]��N	�ye�����^�(��(�O�%�-�L��ƩjG���QK�Dq{$r�+a��x��9\��4�}��*jD
t��m����Z�
U�Wؐ.kܬk�Ӵy<o)D�?�����KQEϷ��bN���nBl��b��5?6�k�3�j��|���n��189�=_�J���UV|*b�0>��˃R�Ū��E`�<��'Y��ɏCi�]�2� (x=%D}n���C�}���
_��Nט�G���њ3� �������tu�j(�@3]Ը��">�F��!`�@��m��}+ǩ� E��?���g�Ŏ �W� �c˖�3�^��"6�%ڋ�T��;�U��d�h{��>�����6��K�X?�$"�����ʮ�����B��=�o�-@�H�6����#ԮR�� �u5z�	��O�9u����ӲF�r���o�6��� p|�c��e���9�;Q�8�f��kx�:)�g]pXf��6�S<�ۓ����$��4jf�N�p�N�TIkn���r���ST��WN�k����4i�S�`8�px��X
W�Q V��r��ڔã���b^0E����,x%jL�NӸs��u^�3[ERх�\'����6��W���A��?`c5�T����B��~4IO�%T�^� ��GY0+������žw��f��+��=���/�YĖZ�	y=��~{���N���a�n�J��w�d��)p9���b���Ѡ�M#c�;a�nH�Fx��p�Q����b��ن�=^��
*q��5���R�e&CT���û����m?���<�p����u��|��pK��aFX�Ɣ�'�g0���0�T7K94�jD�Ȯ=��^��̯*8�Po�+5�֠֐ft��W1*<�����e�[��ˁ�����C�^ƺ��������	�}�rƐ�ق�,7�&9��n��e�O	�$�%-@��H!�{�I��_u���6�IY�9±���ѼUȥR"f�˛[}A.l�/�џ��k"�s�l[ح�y�0Aq�np�� /0sU���_
��Y~�S�sqG�L��H��\y08���WP������p�)�_�g�[�x<={K�7��4�m{���%l �n�|��O��ǣ�ə�B]�3l��ϛ��I9Y���85x����^8�|��^���/������רW����˯{|�0��`d_6�bV�!9�R�'m��*o C�FOԾ��������
�a=�3��he�m�mt��Ay�ɏƑH��'��D:�:�4�gZ-�Z=����bMu`��$;���j�_�k�k�w��:�����*�Q��'�t�͢ƻxe��3�#����$���^�^5�OBh�;�~�.�8�v���h�k᜻�<Pm�V�"�5�@��)��)Dq�39��`����êO�Ihv�G�&��e��Q�W����8�w�dHsi0a[��F����R˰3W}Gl�]q���n�V��2�M����J�KVىv�Ė�5�8� �uKTx��M� �bHCYph�s���P5Ui]����0iekdF�v��"ӈ����'	��2&�O�6?]��}px��� �r��m#%��QSBے�8�ah��RPI��P܎��s�fE-�tg����Ft@�x5 ڮS���O�]�b��:����Ey�7��:��ku��k�걡Q�.H��G�BJ5TJg��U�a�[���r7$�x�r��~9�Ԣ���h�2�����o�z��0)�"]
=Pi=�G��H��Zl��N9�'ie�>���4�ˑ8Ri�
yH6ޗ�[��_��"��9y�"\��H���<�Qpƶ�+�T�N9h������(U�>8~�0 �(լ[i�h�<V�4�$}T&)'L�*���%�wVT����� ��V�[c�Ep�^��-K��ƃK�!���<oV=!�0��	e�Q^�C��S���L�n�Ҙ��u��7���q?!�σ����/�����)y��_Ү{�q���Ú�۴�_^�����Ġ�Ii�]D���D�Ґ3A[��4Z��]ORȺGD�Cl]�"����]/nao�B�rc����a@���~�r#S%�,y��kƽ�8�5^hhs`�jha�Uj�)�}5�F8�G���?��&*�����Y�H`}��x@�K!,#/( �]pE��p� :�>��dN���S�������2�D���IU�,�J�K����_	U8_�^(:�³��ťt���
,bx(���ظ"7"_Kp�:���;{����O'S��[�Z��5�N�bd�;ӕ�eS<ɳy����A�*,�` 5v�=�)}��B��g�
q�,����w�2��K�y"Ȅ]�L5(e�d��Ij��[#*t�L%m��cٞ�QC���Y*t`��@yS{4Z�b�Y-Z9ZNVl�)t���B-R�����﨎�u@���Y�H�ҡ(�yݴw4���gR ��L��1(H�"!�p`�˨
d�1#%�h	�x��?��T~�UV����ʗ;�'�qO��D\����0�⨱�~f]�L4Y�v?8�ߓ��d�7w���?S�$C������6��|����xvdm�H&�R]�_������M�;Z�K;^fs��Y�M�֮�=�z���~���Sd���|%����1㦜P�.Cc/�쩿ߙ$�G�b�Y�]ƅ��
<�k�q�&��˝�˖P
3��Xܛ�Q<���x�-�a�S��2p�w��Jz�61w<V�����蒡K"�O�+Y/�r#�0$��7@���ax��JF^�mM��Z�lcd�\jY��`~�i%�or
~�¥��b���D�������-k���w�??E�H7"nRc�}�$�pON�Q��2t�_qm�Oqu>H��bYcT�@�aԔ4� #cw��4yWc"�+ҕ���o6��"�ش0�kev��@�7����+�RM1���C䁅@r�[o`���=y��S�������ͫ�8�;�d03�Z�����ƹ���w�y����_@UJ�J��QN �5�.nG�o�=�Xیܳ�+�n$.$TԿ7v%^ԗ,����p:"`:2�)��3������U�9�;"��ޝ�&!K��9�;h� ���K�|r9�*�X/p$��;z'6��&WOt�@X4���֠��UCNy*���W5M�� RU����c�i,��t<�܌U��t�?�n�ص�����zG��)yb}�__n�p���K�3�®r�O[Ff��B�I���P��LѪ�0�<�~f������sW�X���-��`�j�ԼVr��4jG�IT;���\���`CE!����瓓����;��dT�+�s!�z�Cw$����`	�3���d�Xޒ��k�t��hr.�P���qm���,���7��G���|]P��[~2��|k�qP���-q�������<b3�y�o38�=�2�H�	�ː��!F�#��x^B^#�1�h��4;�7s�H[X�H����߫��~�m�3SB�q�=�Rן}L�:+K�w߱y�̋��*
�)��%���vɔD�t�'�6�v�Ƈ\ʵO�z1 2M�A\��w�S��w��,[Ί��4ZyN��s��ZZz�&9E��a}iozҤigK'aw��;��bvq���!�n�e�����4j�"���Ʃ�[!'m��(�����,��9
W����S�l��9�%	>��%�PtH�@�� VH���u�*��݊�{	XJ�ȩ�:zsp��bz����X��ZSfd�xmn�	/f���/ �i�(쏗�&�^n%E����25j��oёE�2�C�o��$� �c+i�	�����Ϝ ��(���#��������0\�f�DQ��.����v&�ꆲ_�Kq��F��5	��	���HL�3�$�ό�y�T�zI3-JW�<7y�}����Q�^��bo�;<��Px�֌$��Q}�\��K��[Xr��f$�Xcy&�0B6�w~��e�VgH=� A��w�M<��,��������E��n.<\Q�����*�Fh���)����o�F����T�%���ԧ��bL]��d~���ח�)�7�����}&��>Є�*���x�����������tFf�8�A��T�wY^<s�a"-�.�BG�����[]�YZ(����B��Kg^���=�_a�~��1g��!3�����xp�mkiJF,p�G�o��b:�n�h��6�X��ej54B6
~4{V�& ���"Z-`1���ڈ{�HZ�Үgw3tJx"8����X�?���6�Vx,J�1T2q�FBLp�W_g��6匫ϱ���P������o}�<�{��P�M��k+^�����SE���Z�r�ɱo�F�\�u�T���Q#�1�`��΅g��Rp�驌�j?�ITk������>:8�R���NI�'�/�G�CY�ӲD�Tr柾vW�n�x�e돗,6rOv'�w�������;�4"?���K�V�];��=W������;�1�:����,6/H�Rã��~f���D�$������X�-��P����{���~d�O�kir�u��[5)�&\N�~��<�B��p��6��������%WD�+n�K�(;�	����9�d� ]��
ZMF!�Ly>���J���'H��o�_�gK���NU�TŹۄ}��Ͻ:!G��Ұ�R�Qfޤ��Aˉ�q�x����G��-iN1D!��)LI_R�w�-y^ir���]��[�{f˂ [����R�({9�HY��z� ��M�Ć�����1Iڤ���������|�Nt�gaD��7K������w�&���;�>�ϸ���ν�k�͠嵄���1ғV(D��
5���j�F���/|����M�(]9�����?�褔��m��m��5�����KW7o�p\D��4EU8��e�Κ!-���Q/�9S1u���4���%_���o[閞�����rx� �¶ƥ��fԩ����}3���^��^�|i� �"��vg�-{'�h��7N��'Sx����+����g�n����CH�I��-�cƯ	1�������h��lQ�b%E?����FbÏ�t}&�}r��ƿP� b �.����gc�-_2`KI~�$��ި��{�1rt�-ϊ��s�⥢��jL�T�W��%�0���&O/[��� ^��*E�����1�����U����5?��)SG�M^VtV��u�^����_�f�{�����~�"�J�x����O�R�����ךڿG${�Zr8�T�w\_du��/wFX��iC.�}b�88�d0d�M��y�����.~֍s�*��y����B0H���\����-��蚮��:h ��0�]w�C���6����	��N�ww�`���u?����W���k��ڻj�S����3��ػi�cԛ� �\�i� g`e�Z��`_��'`*�Ɵ��kOP���q�j�;R��q���gr�h��e����w����r�B����Ƅ1Yg���QQ�7l�oRDH�:E����	��}�oy�\~�8b�x�Z�h+�T�Wv��W��W���@�h��5\�EŅd>�����|J��ҿ2[�k5�j̨�$�֔y.L�9�*���~��i\[�z�2,�Q�R����r�O�Y$��ޝ��C�B��������������j�\�_�a��{80l���6��ܢZ��H�^-��?g�"��6d��8��x�b"�]��TS��� ��CG(�&�P�SRz�"�Rf�}��s-�8��V�Ŏm���bJ��F�.���UǯO����8r�N�h�HJ�y�Py���+3�}j��0 9TN��-���k�$oLqqF�L2s�:��.�֙�4l���s$�
�M��	�A6#Ԁ��39;<��9Q��0'�m� �Ž�u�m��v�}��-6mf�?.�m���L�)&�u9����Y��
���&�!�e�"�Ì��S���L�[v�o㬚�<7.[���3��{�`����a�z���X��a��?61���#�e��A�Я����W�:�~�7w�❟{�>�h��3qo9/�r�����ϛ�'K�36���N�2ױn)erHYu�~('^��S>;)�Gĳ�������%Bi�kr��h���+�ݰ�I����S�	���F������5���	�~�bM��i��>Ξ� �����7��"\ ^�H�ZL�t�\�bF_�X��N
��*2���}��)ˣ�����1xCT�����k�$d0��fMXT\�/`^�兼��� Mb�I�_^�и��H�6I�_�G�����g���y��8�׷�B���m��D$3���$��`������#��E�ˌ%�"��D��D��&=���:��vJ�\[�S���wj����q�O��j��)p��w��f# &9[Y=����݆*��n�P��j�)Yq*����@�b �@���~�ig����6���TT� $��N�^��|Y#��_��ۺf���d�aĩn��R-[s��rM>mzj���|aU�6}�F���h�2,�7`� �šV���J�D�(�����]CFEQi$�x^��6]��������t�Ja�?�',����W�X��,�Z,.ˌ����E?�}Ü$H���UO�TKt��%�#���7)�PZ8
�"YZ��GA��9�7F�S��	���,��/ƠVS{sBTr�Szˮ�z�e���}7;}h,�;
n�Z����}���m�S-%��H~M.�$���y2�Bˍ
Q�]�������X����P�'$S	 r����{%_b���jgI�,�ƚ��$o/M�O�#|TW�ϓq��ވ�2vm+�#�c:�@�u�sԞ��="R�|�q����5yW�M��N�U�ux|�gm]��ǦcQ�g�G���l]S�9����_;�I�j��*�f�jse%�qlt��1u�� 3X����N5���t�(_|�O(*(A/ث#�J��ś@M���_?zݟf����O��՞��Y��>��p �3>��jnsw�������l�&�n�BL�gar���IyL�zph;$F< ��]H�ŤOǯ��hC�v�v�ڛ�׽܀>�gY"m��H�_p�P�'V�Z���A�]�;���ߟ����h9Y����F96�7��Qe{\�<�<��؁� 
�Mg'��+���1R���`�R��|��J��%}~p��5j�O�ߋ+�J_�0��5�q��&6C��k
�qm��V"�dx)��f�&���\�R%�wp�0��=xq�,}24�\Q^Κ/H���Z0G�A	���&�J�4A/�㻓Kd�W��*��=Q[�< ��٪Ie�:��QQS= ����2�
\+k=��qW�WeM�ni�@�ܩ����5�C�a����8�#՛��O+���h	��)tG;sxE]���9Ч"��y��1P[u�\�Ԙ*�����t��m�*��7!��H{V�>T�9-�NSG��o��)��G�K�PQs��Re��tyLM����h��.�Ie��)mln��1���JZr�8c`m��((�9[D�����,���O���?�C�2����)�H��Q=E��	?����doz���S3/>��q4����r�|�^`�ؤ��B�(�up���[/��BtB�G2�_�\���O��&��yu�D� ��\*DsJ�
uÈ�������)6��6���5h�i�-*�b:�Q����)�u�E��(����r4<�"DDJ4���G��κ����͇�K�N�п\"��f�Y͞OlY)s�!2�7W;���N���T�%�� J�����v��#a\9�G��`�e�_?_{�I� c�L�n#�4�q`���Ɂ�� ��St���%���c�Q����8u�W]�P�:R�Ⱥ
<��Yn���;�)��ܹJZǇ0��2 hxSS�js�B,F��H�u�ǆ�3o���+p����+|@����3�x���t�!�����a8��:����-����v]��L�G� ��畅��!��3��m<r)l�)�Q�t�I�;���!�T��2zb�5����[g���*�J&���g��-�ZB���{��Z#G�lJ(H[��g~Ƒ���T�x�叽C���7u�����8�а]{Q�Kf�����{����Ǝ�b{����	��� ���@� ��&���� .����6����3�����[���)�%�B�q/��p����EX(�qy�*Vw?��x "e�P�ka0�`v51mE�[�g=���g����[��.F���w%�	Q����N�v�W����}č
��C���v,\_)VP��wZ5GTF�ɋ���Cx����Ref�XpK���bNf~Y'�u�c �"l�/�dѦߑG�=���,���("&����Nӛ_�|#�q@>��]A	n賝~���� ce(� ����}d	�$}����J[�,�.�*�4Z�;m��&Oss���*e��i�C%�]BL����M�Ya�W1HiyPRl��`�Tvb�y�����5(�[���2��O���������3��������^F��z|u,\�>T���(�fWZ[�1�ԛ�օ��,�f]y�T�\]�Vt�*��3>RȢ%A����	�����g�Is��4���� ��(:=�Icm����Ҝ���GG�s����^��]���'z�w�m
݌0�������s����$O^՞*�?�j9.� ���'�;�L�8w�"-�:�@���zh�C/�ޙ�1�=�O[�rs�����,o���x��սt���y�8��Xc�?����4!a����6�D����I����؞W���K$�<��Q���]lM���=�ݩ!v45����V�1�V���L�LgEM��Df�َ����]�O�S�|��z��{?��2��4���'x}ꄥ*e�H�$��s%#,5�p>�{��O"�n~1�F��0���.����u�4Um�ٌ�JPTR=*r���J�r���km���Α�����K��,S�����_�Jϫ����#h�ozd�k|N��Pwe���?y�(�W-�1(t[P��5s���|��H�G�����HH���]4�{�ܦ%���V��8e+*��1���W�fm��ky�>��}:ё�������Ǯ���;?�^��Qb�"!?�\g�䙉bh,z咠��t�ѱ<!A����p��f��b=#��6u.ʨ:���"�mD�H��m}��[�3y㋤�'B����^l�7��������Q��8��}Q�*��eK��h�G��r^^�u�(t))�4���P�e�;><#}��tj�p3Ҟ�o����Y�6�d�2*�`9�,���:�7�C�77!�f����Ý$�`���mj�n7�TN�ؼ ?��e�l�x
��/����E�<�њ�g�3��t����@'��Y�r[UŢ� ��RM���Ɩ�����@��}!QI�Iv�����d��R���{޵6+�UC�YZ�+Ѿ�&5'�ϟhWʓޕ����W����-�����U3��\��V8�'9�G�'~�b�u)}�|���K�=�S�յ�"$�Tx?������#�qp[��t�c*m~��D5�C�o{f�7��%
�ߥ� N:�H�p,�aP�ܸ=�1#��{+�J���;
r2�]uQ%-�6�l�OU�ގ��z���$[�e�(�� � �b�%��C�T����T�zl?S3u�9�����:�ɮ1���&�C)Xvb��Si��E�M]X^���4$&D=�յ@��<���U����Jף�����A�e??
8�G�K[�U=�nl���"�ʁ���Y�=�]���h�ᑶ_FG�߭��S�u�"y%q�,Ւ��5���������!�I ��ַ��#~v��WZ\*a3%��_o�Xގ�g]��c('��ٗ���]�	c�)^���Byu1f�3k�|�����Z�n�%�tl�� 7��D|�d������!_��U)^{]�冧T�e���4I�J�k�4$���#T���"�M�;�PHp}�XX�}���g�3ĉ�S QAA��Jd�MΗD����<ɿ�ȓ�K<a�>��k�7A��Ҡ�ǷԂ��!]��;m��Aj��sWA�j	��]�O��]���3M�����P��1��I�{Jȏ�~5�]VK�x�#�B��M蔓��jH��v�j�_��E
d�n���o7��O�5!K/�ӟ�?�<�0ld��>�M.�Z<.�BQ�֖y��as;7-��d�K���C�	�t��j*���%����4ˌ7�S����ߌ�@�f��� se�uSӣ�V��N�}��$j���)�����]f.��x_@Yä:�U���qֶj} t�����Mֲ�Q�#�P����,�j��6�C�tVI����S���?��>R�Ɋ��+4�Dɞ�1�=%���<��ф�'����gi�(�]�F��w�!`~��2�f7��US���������a 2����>k��0�>d�/hp.���2�,�f�i��8 3���q�	 �)��유V��²���uK���������ߝ��-*k��Lt��_ls9H&Y"$�L�ZP&p9w5`�|O�B�(��"�૊�����ɷ1��M�����zQ�h<��W�Q�[��.=Ꚍ�TX�_[�����{��u�(;|����B|Rk�t���bx�PU��HI#���C�~�ަ/�s5&�6��e&f��o|^XnqCF�����Is�N1�r��":5]�{ט��,X/0M6THV����Җ'N�7�� oЗ�-z�8Ge��ޡ�ͽ��l��J�u�*�3�W�^�ۺY�������ߴ���� r(/��U)�^��&�N3�@Ԓ i[b���p�`V*�ӫ�L��C�N!�'5�'�%+�P� ���k��7۱�!��n.+
YӲ��q�M��;~��-�E�?�K���[(������A4e����m?L����Z�,��4PM&I���m^^��hRK�ѿ�������"��u���e3��2��q��T�a�����%Ơ���~�����1��b\����ᔒ{�Mp�¯ȴ崣�.8Q��<�x�?I��w`�NAxH5�t�t�7�
��R[�D]�$u�/�6���VP���ef��Uꚥ��#򓑢����bH:GXJ�X��5愃�+��yT�z6�?b�Q-k]�wr���D"�8α��&L��0i<��H�c>㠌��K�a��*�6L�!c{\��28L�򘫢֯�3�H�j����!"�qX����)@ 9
c9��|�d��zw��6���WN��7���UdW�y��Ȝ[��˟yb����CZ���D#�K���⎦fc���,��� ����gm�Y0X�S�k��@�1����?CYhb��>$���q�%K9�!����]Q��P�~�x���[f��%�҄q��l@b�R	���z���'
���*P4���w<.�Z'�j�@)lJ<��a��*:g$�Q��*�L�c:�	��r�*�_W�$�тarFg�F�3��t�s$�7�X�C2��v�X�)��G�ExL��Vs8NZ-p�]��¯x)�3�!ED��P�N��mr6��*Գorg�gGr,U�;�*�ىb�zO�QE�7@Fw+a���R��n�ٗL�l;(��K��A ).C��WM�W~w�����7,I����ȯ[�������o.�&�1�F�ٟ� �����&P}E�?���17��(߃�,"-��y#�O��˃�gS�b� ���-�Zǡ�;�nX�1s�_�"w��t�hv���h���܋�k���7���oj5�����A~�J@���ȸ��Ps%���w�>o��Kz8��&6p~��fD �X�T�'~�,�ޏ�-�S%��̊��Y��;��>7���nܗb6�U�q�ZԢ�����:j
�1?|`�[c��Ur��]m�V5y���~�1���rn��c��VnC�sV���xF��|xҧ��fh��!��`�����4�����Y�Z��0#JEM����˫xmh ��׫-��?��$�Dn�W(ik��}%A�J������rk�r��;V�TO��YUP!(_/�)��U'�M�#�˺�@���]J%�[7�Pb���9箥�7%��3>"9I�ƥk������ϿxC���+���t;(��`��!n���g7�g�O6̒IF� Q��dẁ��ѳ}�T�ȥ��
���j�1l�%m���ٽ��=�fF��F�ں���="�Vj�4�G~Hi��ۮ�RC�a�?h�1��z+���O  ؠ��g��I��f��[�ʋNL��#
�'���o���N�s�
M�z�BaY	>�6~�,�����c�y�h�(�z0Jl�+)�O�5$��_l���"������¸Ԁ���/&�#)w,+WRT\/l��ހ�]��k6PƐ���@x\@�!�[�&s�o�\3g�?�yߕ{DI"�e��M��G��a7��$���\1O�faZp�%(D&�����n����I,,�e=�7:\I�\3��T��,q
pv<�f���q��A��B�9�N��y^Ixs��F�<��V@�1CT3�����)u�k�o��0>9�JSH�	�u)����Խ֧C����,�X�ǲ�t��B��#1��,�W(Ƙґ���&��|�{6�H��g���q�%x��iB�q�hG��6J�N�G��py�_����a��$7�n"��0��s��*��X.:4�x{�G����c���П��o�el6���;�
��R�v{����ۛ��8.'��p �8tѬ
j��xp�>�*����B3�qz�:素�,�"<)r�{ʼ)���?��e���-S~����k��Ӟ-k�
>�cVօ��}Z�hK������T��C�
��MW*�`���J �������U�4��67)���1��i�1*X\6����\��1@�G8l���ª���Ὁ��)��\�SJ�3iW���Ji7����Z��A���l.
��x�}g/,5!�&	0��\j4<�~;��#���&���w��US3�8������Ɋ5�oT)�U�eB{iO���VZA��{�uc�p�by<�ĸ������aPt�	���8
�J	��[wm|eM��寷�nZ�K���q�o'yW
����Gn�6l�rp�ew���@p���lܾ�/�]�kb�. ���q�Q쌐;��"��jY9�Jў;8�+5�s)��="s'�m2a���_K���8��DC��t�Bj`�Z����;��Z� ��(Q���?ѭ�!k"�Cf�eܺ�J�s�����6�	�IcbǗ0VF)8����C�� 2Y��)�jd�&2�&Q��g��U��3����HIеw�,�\�NK@�侘4��7�c~���~M��t���{�k&��oR�Υ���*�*��ɽ <!N�r�Zӛ�t�!�2���e�g����hj�T���瞔�KI�߁��j;����Щ�;�i�(zo��X��4�*�w6��Vi��	GNo�
��� ��o	cӐKyЖϨ(��5���`qJ��PK/B�l�_�������ܕZ]��Qh�Hz]��ۛ��(���y�?}��\��x�h�ņ�S!����BK/F�0H%>GN�uח�O��H����O��}��S>o����D�+�9�<>n4�n��w�`��t�\x�C��*w��}C
�������̳���M������|���w�2��L���6� 	u��czf���5��|p���������Ф�����w�m�6:F��=#�`L4���� �y�ݴA8�:!8��l;�1���4���A��ű~���G0���Ǟ-$垗!=�7��Y�#$�H�mW�]����96*��j�����w�>�䫰(�c�)��,7�y�_U���[��wq.m_(/��Y�ɛ=O+dJ��s��Ѻe�d�2�����C��1vR�b� fe|��-��5��&�m�x�`����?d��ݼ�_|m�����D�d_{1z�]���h�[�n1�x�L��Ƶ�i�t3�M�1|R�$���!�{ۡ���~}�ǃ��6
�D��G�P��-"A<|M��f�?�}�/Ds�u��G�ش��c��%Nb@��>�P3�N��3�c	������K�=�&gm���`�".�ǌ&��حahq��P�z���aսC��i$-�{s��Fq�<6&T׎��Ç�R�_OU�	G|�ɢ�9|S�Lp8Bܾ�D!;X���zMJN�  �喝~�V�~���t1��$V�A���L�S�w/�G��&g�
�A��Mp�l9�g����	��J22���5�8^
e�"�n��t'���
%��wq�6(�|�*d���A���}9��`㲤��|q|���]쎘���p�>���RbX��t}(�"���wh�#7� 0���`f�"@Cd�dU�'�U��aJ���܅\�&\5����/�^���_X��mejv���<>6���u�k�v�'$��Nx;jv�k�3���S�*ZU[�y{�[r"��GO`E;s�D.Q/����?&���u��z���*�k���V�rL�h��&D;"O��j�2S^���ϨQ����K"kr�P#����1U4��[�?��*�)�D���0���M5�P�Q-��W6���B�.�[�R��H�����7+T���nE)s��@�쎕jX���G�x┐��m�R��.:��0V�u�����o�"}|���D[�i�D�����k㲂������ �+*Z;���>An$0'N1�e�����"��͖"�w�����$���*>  �8�C��2@��yb�*8���RU����m]�-h���):��3�@��^� B���f�-�F��_���+�(n�V�����&��F��4������B�@��I~C��F�!����S�����@����h7��.�D �`>��&�8�Xb���&}��Z"�>�54����Jͬ�/CԂLG���BX.M������^�,���q�Uh���'=	�h�T��%������/9�.?NE_{����hr*/��{�E"��{V&ykL?<�6u�\�uժo��X��͗�Ry�;X1l��Q�t%�sC��
�?����[��A��Q�90�S��<����e���G�]�׭�Fζ6v�����UUB��+��Ȕ'/]�6ߥt���[��*I+��0v�y��!��[���rSch�YX7��Bp<3/�(�3�
/H�Z�c)���<81�N^�܃�6�DS?ng��P3�P*��i2�i@� ��/f@<��g��LЖ���/���5�h�+?�>	����s���ن�@��\p��Du��W�T���*n������O�|�ϵ0�	�O'Z��U�#����D���V��B5�z����W%����]��}B�&��ƺTQV��o[����i܇l^�'�^m@����� L�,eY�D�d߿�:c�?TК"�f���N

~�$���vI������^�G	�Ko��6G

�3�d��S��&~m���)|\f:<��6�FM������>ڠʍ��%�J)6��W�0������0��Wj����n����	�����t�.Ǵ}k��P�W������˳��O�����=y�4��x{�y��BN���s�=EAO�к��ꀫ���v�E������~��;�p��c�?�Yz�-kN�dpv0�f�����?�Aw�*��w�n�d,Si����dO�n�i�7��-ێv��Ah9��Ŋ�����y�RӮe|� )o�YmV���~�/Xі�#���NϿ�3��Z��$[(��[�&ڔ��ފ���k� D��w,&nGA�hi����Ar_�hFi/�1�\#���񔁡�k0�clx$�����g��^�U$�f�/^��: �D���\�w8z��(	����Q�xԩ�`�2ѧ]|�(�9�ۘ#'�7*m�o�5��%7j��o�����"78rR^ⲍ�����Q'��w�'��7�#䓒�9�]�����G�4^2��q�%8eU���q^����;�|4`�	�(�LU;W�L���q�i�[� � ���-d�g:�}�-�,�[��J����3��'��θ����UG�,���u���A��H]��A�l�0�L�m�]
�%�ޟ7ĭ�%xc�?t����KI�eq����/�ڭJm��]=3d�9}�z�hʫ(m���P!�d����1C1'���Hr��L$;x������l�G(&���Æ?O�i���{�}��9X"&Zk��^ug��]b;�%9�H��!���^�Xm��t%}�����Ce�~g%�s�758�W$���4|8���*�l������O�.�b�,
�+s:��P��1uH���^.�p:�mA�ء�,����W!�-��Ia$+�Kr�z��6�� �}�"�E����t��ZgW��I�y�P�i����z��� p��>��Mqʵ�kI�gg���H�Fz7��VxZ���_'��3*a�͠J�K�=�n���<K�}���P���
[�+�L�T��+��5H�faE� B���9Vo(Ο�\���ZSS߭?(h�jƮ�zb���Q���m����_��}#kb�B���XFm�|���m䒒N"y-~�����Չ~��|ϔ�GL�1�6���M��	C$��v Y���JB�E�h�ba���/�r�#3�/<�pB��+|PGZ�z8��>�#R	�l��Q`ëD`������01e���>(rA7�']�W�㞊(쀯A�Ɲ�����<��~���-��EypO1�ɚ}�s�ɤG�މ_2�л{
-�_J��

,i�C�c'�Z��ֺ�]ܦ{�N)�lj��Yd�"�r4�l��t��K�x��6��v�O��&�ǵN����Һ<c��m|?B����A�t���%Z��nv�=�%5����M�0�ʼ�����?��@f�Ц'�2�Yl�0��D����)�1>� �VӬW�����v8��F�x�L^��&�v��=�>+�6��b�7��S��n�}RF:����X��R~�m��˻���{�K�;��S ��2���� �V�7X�xJE�UC��q`��#�x�Y���ۑj��&�h˦!����G�=���;h�V�M��Hۣ+������:'�,).2����w�ճm��+�E��u9�h�*?.z����F��R3	���ա��&����L�(����@��|�����/�.��{� ӊf䅊��f�>���E�a�~"���_�V���$�^�'�q9�[�[��?~ʷ�T���~>���#1}��f�M_���3�ɗ�T���~O�4(���>9x������_a[}1�պ\ba���i_H���<��=��'k�qZP	�5�|�KǠ19�rH�j�{�t�Ka�?g�'�����(��
A!��Q������d>�ъ;����Nq��q�z^�wOERi�j
+J�B�033�2TJ�)�)	 ���P!~,�p�rK�,��zv��W���R��Er� /f0������K�X���oNc���Y-)�&�j�$�,x�]�ٰ:���oG�PG�z�&��/K���E����۴���b.d�i�&��	�o�ǎ9Z�k�Ŵ��fW���?���z�M��)]�@�����x�?&�Yc�R�@���v+y4Ŧ�&0]uB�'��pO����[0K��V���8��IiT�.A� -�g?ԫvk��L� �DR����$#�Ӂ�O-lL(��Wi�~A��ۮ�	3�-Vik]y��ƦhF�M�-��G��^�2��钮��i�wS��$!&�?���2\�jf��.���a����׼%-~^D�â���:��X�ho*�W5X�ǝ�H�E�C��oS�ȅ��(Sf06�����8��+��c��0��y�Z����\��pPV��A��*Ƕ�Ui��=�p�����Fy�u��gdB�..>�m�r��&RFљ�����G�e����}sk�q7z�o4L����A���UF�<�����B�Kޘ�3(�����j�b�o�I�S�@��
�)Iq/(�f��~��Z�|7���B��ې]N���>K��&�5�$�m$��4��u���෸�|f��-��Zd����bk�T�T���u�8UG��g�P�;�m�Z [HQ��b���Y�A)�\�T�)��4o�|����-I�������q����'����o엂`���W�φ��y'�?k* �IF�{�\�����*A���̤!�V����Mo\�9>�"kɧ}����u�-x1��`$���wJ���(
�ᥘ �2�|���d:�*<���4v�C]�Q��Qŋ�"v9��Z������4�5F�l��L��p���unR {� ¿ߺ~rIr4�D/5���%=��k~��
�/;9
��|w�E*��S��[ܠU�;�92���w;D�����ZvBs8�6{>_�� �3���d-�N�[��	%��RH��&�/d*�I��h�m1|�����(]�������*϶������\�P�Ar�_Q�$�&��dyu�ռ�zk�:s�H
�fA/��4(0';�ri�ٷ]��v��*�BV<�K�[W�.�^b�l�H`�H��&	u "�M	��O�����#湶�[�D��A���i5V������.}R��''��A�x2~��F�o ��b[���/^O#,#A˱μ�������?<�-��QFbq1�B� ��5�����;P��Jw��=8��|�6��쌱>&�ޟ�ܷ�IK�Q�}��v�๵0�rP�_t64�=x��cZ$��B�&�A�.<�N�H�Q�RP�
F�F�ַ�h���o�I�<��u ��cT��� �jV9w������+��q��_�N��.�Q�{�{��+��{���C)X�f�����tE��VO`���uL�p�B�!�.b��N���-q *�^�ݺU'nX	v� �!���\)i��<�l(���p��b ���*��(U����	e������-���D�O���.��-���"�C�,Rp�}q����y�'�'gB�M�ش�(��IVW
��xz�<�-�n--�+{��M!�Z�m���J��Eϔ0�3cJΒy.�
QSf6���h�����=��������4�r�]Z�).v�9b��p��9h<�LI�
�v�O�0�ꍼ����
��{��x�Qa���#�wZOL[|k��n��{�V�D �j��;,���L��Y������=O�HJ?������UV����Ӑ����#��m!�G�:ie�q%�\�y ��y���1�=�'��r��+t�P+ɭޜWPډ*��&x���,��X����69(8Α(&�!�{ꮬj�j�m�V��W�]h�W�B����9#N�e;�*�T��)n�\<�N,rj{VyX "�G�[p�$A�[@u��z�{�\	�� ��d}��ʷ8�xAm�����:�E�4�}��&��#��y��p��MMу$D/�jV�$��A����/o��>�.
��n���La�K�8���a�R^����nߋc�K��0��X��$��#~MϋtY�E�x	�T*�i[�����p��� d_��\�R�N歈����u��姢�'y~��y��{i�=D.�C
�)t��{j(�TH]�.n�gNT����1Y7l���:��XHP��ٻ�o7#&R{X�,�LG�ATO?ሻ����n�� "�`3 . 3}G�	����R��h�曗���y�Z�-��Q�z@���=���; ����G�	<���%���Ål�s4<M�@�v����҃��&�����w��E�����T�N6����1՚,SZ]��؀���е���Ό�&"]�t�����5-Ė4S��i�li���4��->��%��cD��/����LE}��N�ch�.c��bh��#>����t�����?��� 0�y�ъ�<��!��|�f��4;t�F��DX�3���t"���0�I�M�Zb�1=�7珸�+�Q��铮��b �$[�d��=��g��Lzm�đ��J�'��z��߬s$������t�N�e��@Ve��/TY4�(rs����ZG3������g�^�1	0������p�C�]��C�U�Vq tB��uF^`��p������W!W3�����dR�N\��B�>�
�O�P��{�{맪��!r7������Ke��_�W� /)�1�% S�a+0������#���]������f^��md ƽ���1)���5E����o��j���c+,|~Q�O'(a�������8�6�¥��L���=�ݪ�y�[]�Б#⵷2Tc��O��|x'���ȡ����9@�e��%ZB5��w�4�	���=W|/��)5Oѥ���'&��w����-|�ɜ[dP�n�{��F�Ĥʢ�-ϢѠ�k�B�uk���{�a�s�׹��>��?-���Ǯ��N(�zu"�,�0j�Bͭ�]��Xz�ȍ/�}H��[�§���_�f�C��XMs��ߟd�~+����M˯Do�4��)J^�S��jţ51�{h� ˪Sˤ�;������ԥ�6)J�-���f�Q\�E�:~N��*T��sI#�K�n#r谝��>�2p��τrr�����<e<�����Q����Q�^�6̦���AZ�d��w�j���o��t���%��l���$+}�e�F@��ۥ-|p藕�Hݽ{馳�$W�̰A�����9��pɢA��a�����ܽ/������v�`�&V5�|�.��URms�BaB�<Mo�%�������.�#{�V��P̱���g�l�7�ܿ9�a�Ϯ�2��7.G�;�9�*�U��?��0�GV�%���犈d�Cl�J��3t�ѾS�lK�e���)��?�!@S��=�z^4��	����MRl ���C��� [�9911�U�����q��(uXlU����w���"[�M!	1�|�7e�ۊ:lk��4��-���߸l�d2�	�14;y��X���������I0��&	q�\���x��J	�0K�_異��������Q�G]}x���h��]��Fi��@g��=���؄��eRo6�)��%󹚪�����3��ƻ<��7Z=)�f�����R�8V�HE��)v�Ժ �
��ۮ&�g�������6)�1í���|���h���i�Rc6G��O�YO���	�.0������̀�Y��W�	Q��(4��']��|l|�ѭ,�V��T]�a<]`�9�<b��Y�}p�Ϊ�e�_����;m�gOȀ��ތP�Ũ���39&���/C�Z����gHE'�	㙂'xS\ͯǾ��A]\@�����QА`<����9P���\`���w�j�(ѡ��d�M�nA���..txY�p�N0�}֐��:���h����������.�K �� !�$8ww�!��������;�s�=w����Z���ꓮ�����[�|�����:4_w0�uzz�����M?,�l���*$�̭�Ժ$�Kx���s �a�B�G���E�_{u�ă�-2��t��7�<�X��X2�H^���4�B8�r%��ǩ5k��i-�05�
A��������������fJ��FZ�O�#HŶ��ĉ$B[}�6[��ĩA��R�ڊ��߉��<x��]k�k���O�;?��X5��/����� E���6v j��f�^�l��b�'�?���t�V�GbP{g�yB��RiD�(��8�xs�j�PE\�"�&4|��
i�
`�ݿ3 ��oK�W�Oĵ��Cz�qRv��Yc[*���U���tm�ޝ�6���Dv����D%jȒ�8�sM`������Db���;*_RIf���0��6�6*����URZ#���hQ[FE�$��?�q6�5�8�ei�,YQߠ�fO��� ��ijR/��z3vi0y^Pl?�O����x('�-?����¥<M�N �0�*�9Nk��3Fc*f`���/��I��O5*9�k����pz~{ι��5���G;�{�~�΋��^�V�t�S�P��xƄ#�k,5|~+ ����e}�{��}^�V����5��|¶���)��Z�j���&���)����Ο�IȗZ� �k��_��&��x ��$���I{{}��Hx8��">�ࣾA,�������P�A��0�}����q+r����^�]6����?�$�s&~�����c��f�SO�����e�TO7��5v3K݅��	�b���G8��Iv7��_���a������?��e�X�r��=~m��<g�1�RsL���*���{�i4;f|t¸�����(A�U����mͫE����ڟnW_I�Ee�\cO�z�����91�.6h�<�
A>�\R�SyH�OJq6*H���xYj�_�B���[-ޢȵ~ ��5a�ջ�p+0KӇU�nt�?T5�����	N՘X���p}_p%+M9�(��>aʔȂ#�g'��������<!��	Cq���^� AUuYh9�j�jG���By�s�ȇ,0��|�4<�@Dz������)O� ]C"�oA�Bi`5^�<j�����a���+�3J�ѫx��<u5�_��m�A��� ���A<f�d���O=a7����T�������+4Ϭ:ݦ�����L8���a���nb4�p���љ��d&�J�I��G�і"�ţ��p�_3���|���A��.w�;xJ�°���|p��{�:	��1�<@�e���
��� ����������&\x�%�G�����B��q�Î�pˢ`l���@��O�8d�Ob;=$jt��֝��Q�, ����E$h�b���9���fb�Iv�\r�8"ŋ��H4�x��p#�R}n���7;�	�W�7H�T��p�H?�އ�Ou���}�� @�lu;���(s)	��Q����6?��ġ��1�ʅ��,B�A?RF������\lǫ�Fi#�� ��o�D:`�We�4<D��iB�J�0
��[i�S����Y;�lJpJ��>l4���"&�C��ב}��CB�NF�j.P��P���.������#�唞ܱ���7�� ~_� &�t�|���Gh��VoC5��U
��P-��������YR�ѩ��/��
��|O��E�������v��,�z��w�V���j}��
�]�O�+�߭�p^.���G������?����M���%q[+�tëq���\��_V��*�������ݎ}���:�-3�{���J�T�={������Ɂ�9�5�7<tD,QS+��
�6�0�8�����D��2�wV9L��Iv����l�.�����Lu-��.�u�R�i���'�w$����i��<�+�����]ቻ�=�Xy���8N�p0�<ɲ���ܾ�lk��v��f���3^�*��}0�C6/d~@��������S�pn6��=|>U��ge�_i�ƁIFnH_���!rY��Yꦺa��^�a�,���X���IZѸ����AO���HΆgG�/pG)v��ג���69X�]ݷP�.f򔠷 �E�wXk��ݾ�x��K�. �5~S��@6'�
����~ē� '� oS���"�q�4F1Wh�ʪ	q�S���u+jT��]�UO�(Yyq>ABX��L�R\�25-�B�Y���2>�}<_������g�!�k�3���D�j;])q�7�[���8ӗ^�<��6�`86|���N�$�Y�61�I��B��$U���(�o����.��B<�r���E.�?��^�q�ֺQd��XY��ކ��U	�M�{���
Qh5v*�>�B���/�7��{m����_![(�Mb�k�(��}CkD�9��2�l��ݜ,9�y��1L��XF�S<��9FR-�<I7jR��%����Ǘ��F���:����_%F@VK�z���`Fd	X^�Vi�S��G�6�8t��7G�@wM�Y���ֶ��xpl�������0{��g]�N�;�eD�S{���W��~g�pʛ�-ץ�i�rv&@���5�-���u������R��O�l{n�nW2������n�$9�����3qn�8J?�Hm}L��>W��{ Y',Y��G&���xIsZ��V����C?�͎�Q�w@/�ѳ�:����3<�܀}�ݸV�~d�U��B�CA��;B�barΟ��ט#J��ʪ�������-�6?� N��;>M���-"�XQ��2��W]�b�@Wo��ێ��W=�n(���i�#Ζ�����Y̛�Y���o|�Ӡ8R_
Ч��~r5�2
b��́����>�%�UC;��m�Ű��?uʵ��3U�87�8q�0�Os��Y�eM{�����\?@rp	O���z:NW��g̏ԕ��u���yS������:�
�o�&�~�f˪U{#��K�Y���@{��4=��Wq2�]����&n�8:�evb��I��5BU55+�j�\�:��?G	�+]'O����GI�-V>E(V�6:���GE�#�n#�I��φ����Xٷ�	L��,�ԕr1���k����_p9N-0`�݋�4p���.��3��r�"�_`V���D�p�֬3F���$��LdZ�����"�G��/i&B���1���E��W�^�\ߍ�6��Ce��}gH�*ƣ+og"�a��9�qd/�����$ד�_T����Rr	�C��WD�K��yu���/�rAhE���;�O�J���>Zr�.a���Er���;X�f:�4��2�<�-REE����:q�ܜ�e���O�C�pd�8u��슳`	L����̶qw�,5F�q &At&l���7�V�׼��q�^�u#Lx��l5w7DŞ�t�$��qz���ʂ�Qj��x��˔�b��͉�ynjა�׷u�ʋ!������I�ЍB�|zV�s2�n�l�U%�	�s��H�4\"{���4}3r4#��> 9A~M�^�*-�I���^!�g��42�(��t��dE�b����$6��T��% �8�����~������!�'\�	�^ ��Aa0 n�#�H��i X�F���AΧ���KD�Cs(]����%��w�S���o�%-�q�&*�u��Z.�6SH�&��P��R%]� �l�ЋqVq?]с�؅�7��lcC_��,��$��_yz���z��
�̬=u�G<�6�;7��e�ǝ���E㉪��p�����{���ֲwUy;���(�'B��1����P�6����K��dC���:����fV<n��[g�ۓ���2�)���c�5�M��\B714�
��Q�j�PG_����mn�ۘ� �Hy���C~��@r2�` @��Ö�(�i��\�Ւ���'����)2W��%�^�i>�����ݯb��|B�%����=�_<�D1)�8�8x��I�1�ɍ��F�?��h�[7Mz�>�l_#�7��Z^]�����/�%0~*�3/�6�m�L(6¾�J�\�n��KrL�[�Ee5��u���Y휪LV�Z�5ˋ/N�p݌���V���gH���2�g�\�_�&�C�-4�M�T�s��=d9���?+��f\��|���Pyx{��?]фK�P��ɀ(Ah�*�(12�>A��y'�Ʌ%:�-�S�����;�N�!"���8`{��绦�O�Ĥ� ����|���HJ&z�T�>G��<��|�J&'"u#�!�R��j/F�%�����*0(%��z/���Y���xR����.�z�f�٠$i.7�}21�S�D�,��\����
o޸���wՇ��?p��V*/~O��<mqjQ��i������I�V0��VT�5��97h.�|�f�@lg~�����N{�1���\�j��H�=s�ө���q�tFM�@�Y�P
��)D9w?��m���?ؗG8�U�<M~�t	�K�����������K��)I��&j��/�j5>�V���FE](GҰ,'�}�t�b��QS���e���1�?�}�0-����݅A�&���+����b m_olNLv6p%�1$uI��*���{�7N����=�d�_�lKس�v-	@�> 0����q�s���ab��87!:x����Yj��s8�ů&�����i�����R\��9@FVpxȨ$�(�<�F�Vq�֎��~�����%���@�(��9p�#|� ��wC��]�Ѵ*Di��2�%>�|2�ŹńqA�5�[$*���&[� 8R9B��SX�Ê�'$g�O9��1$�ݍ�>���B�����OW((!Zʟ>���nQ��%\0$L��q4I���o�{�2�D0St�'X��
��:���m����.��$1�d��2��vy��A��
%�p���ԗ�W�ȃ��=vwId���F��B3 ֔K�d�z�g���/���Kr��k�Q� !���"U-I:Pk&�R�UAX���]���&%�2��ʒhxDۧ�k���ZX�VG�a�Ƅ	�u�ϲ#�ѯ��؋��j1�[��P�Z�	`<[��� ���8�ܗ��ρ��=��]/pP�?Q�R���,ٶ&��@ڬ������oi��]7�E;���jB�o媇������I��I�x�	��>��SB֋�/j~C	�<([�Z!j󼥲$zi�iǑ'�6L�/r�MAK�x�hV���(�K-B@���׍7;�6R�R={�۽j��Q��/p��`�5��"��MU���	R��0�㕛���%\�/t�*%��N���)CQ^�͹���˔!�
Mq�B��wۄ���F��c���ѧ?�cI�'e�r?,fy�v��"=���gqF-����R˲�H�/``;Ey��������^���?5�pC���z���H�`DÁ@@\��+9B�7��/��
���#���
kE�g�u{-+<�t��r����;1��ѥbv���NXD��*����c��m����C"(��-@Ʌ==,���1`��[R7K��:�}J&�,����1�$W� "� �:L�sؖY?����>��7���g��j�z��b��E�Xu=�r��Dt�#����X�\�"���6�K������B�'m���#��9����,��?fe�zQD����5M���j<��n0�G��4�6O�����G�dj0��)��Q���h�&Z��Ge�wZ\�p<�=v�Q� ��oKO��||o^���n�Z'^V�39�y�e�3�'���C��P�.4�6�����?5Z���d�s�9���,�r�F%B�o��t�j*וh}���`�<����cb���A�ሹG
6���������:߮�m�\=��X�k��.�~,�\�
�j�M�[�M~Q_��6�7��$���e����㺲O OZ�P����~y�5zK:^p��D-C�o[��n߫#arB/�(ֱ�=�?C>2��"d�
fJh�^�X�l8��^�;�������St\� ���SF�58D���=�� �8
}�8Tie�ŷ�QH�M�2ߦ��;��q��A]*F����x�h���I��)T�����!�f�Ǝ��i>���������"�wH��uһ���<�Ќ� a�'g�����tČ��B�E_Q^�0jAeҺ�T�-�$l��)d{�.�?֜H�ڃ�y�s{��o�$~]�������� :9����T�7��J�*�b�f?\,y���-�Qr�D0� �uG��g,W���R�=�mV��m�O�U롙�����g�Vi��c��%����:�v?2o���y��׌���ay��a���+���ɐ��t�V�\vϓ�7��1:�r^���q����бU���]^q�h����ܨ\��R��=6_%��ã� O��<������@(��j�Z����e����0��y�p�;�5�� ��7�(��Ȇ�9K�6��/;�ux�C��wy67��j��Z�_��}��N���ƴ,�o�)c#�BJS7f�����xD�q>��.�QZ��b�{z�}v�!�T*p��HS�b#�wM�����k��7��t��TJM3t�$�����܄�}�6���P#����!a�@QO���M�䕟8�8ո߈�o��|��]��2E�����I�%�B�
�8�=����a-�3�˩�|���In��j��qzd�ihÁRڼɊs8<��=�>#�����}O�W�9����f��,�&<ie�^�t��yu��ٚpz��G)Lv1�j~;&�V$���\c	�lP�$2o�����*���T��g����f]��3P��ޠ:	��md�UY����U�-빩a�tM<���Y	���M�M[��L�y����6��UQm�m��k�(���An;N ���;�;,E`������##����	v}��R��v�U�������È�:�
����&��B�V�<r���[�'�dVs����Eo~ߞ���OqzR��,R���]�U�R'u����U2�I��������ۻG]2k!�?��ր�E'iȴ�v�2m��}�1W��hyb8;4�a�μ
_����_��k~b%��5�s�ޓ��l-&���ro��%~vӡ	B�ݨ��UF�85Դ���+�M�g��s2�}Gs���D4`e�Ĝ?Ww��
	x�E��)�	���@`��d�ֲI�)���4Rp��9:�S��Β��4_���\˨J��C���K�����qi�)�֐C��)Ir�3�Rɐ*:jPԱwm���#�kޞ��\�M4�썷�{O���E; ��e$9�9F�!l�]]���|�O�aXvR���#�^����mq�ْrnj
FX%m����bxkN��
qGQ�*@V+����m�V[�n�B1G���_u���
���g�@���Z�tN��������uu��8�Y��H�S'�q֏���m>)��F�0x��x��Z��|�<)sҨ�m�f;�r�~Dƹ�}�I�ש�u{n�F������[�Jl%c�I�6�KН�_��z�-V���(�d��qG�F��|	�7����,��mP&&/MC	��[!�c(7��!÷e��=�uo��}���#[�[Lj�V�S毙�G�' e�o���W4��5���C�G~��'���->d������M
�������]�f�S�|�LN���c��G�dѩ8]q�[��s�BC���Y�����L�4r�_��|�6����9q��Z��a�w�	�P�A~kC8�>|��p�Q�8cj���Y��QB4�^�՞��H�i��l_� ���[���n�z`��2̑���쫽�J�u<���[A_'H���,D�[]"daj�(;D^u�Cea�c�� ���1��^��nǁ8рi#C�ё���ئW�n�6��D�_�9��*M�i�[C�A���Җ���xqR3���*	mĵ����N3;���i��=Dn��G�W��
�UQ}�rn��(#,҃�)7{�|N�<s1������������B��<w�-�d�y�?�.
A�9�f_� ~��D�_��������<�#-B�}� wY�Qx��nGZڰվ���J����R�?6�流�`?In�y���H;H�>]�$u�(/���+��_\ z鬁��l��:e��Wk���y�ި5���%䇻v�~{��-	����9���H0�3ڤ��p���!2��Q��p�=J��TQ�7�Z���V�'�՞�
wu�_�E�٢�cb�=��!�j������*��,<z�'6��u<|��2_��*�o��J�o/X�W�s6F����G��DI��/(a��T`��Z�Ji�Qv�M�ns�ϲ��,��?m �$ 0�0]�3cȃxW#3��ʠ?���# �}�ж?�`���$��Ș`�*"��{0�l�� #@�"��E�gX����M ��T�e��>��͓��(��G�������jD�uML��T��%6&�NN�T���x��H��x�"��Wƿ裡O�����������@�s��Ռ� ���\ɿ��_���@�E��:��r�r��gD�倱~����b6*"�t4����|�L̍����_���'��ؼ��I�Þ���IH�L]�7!ru[�/�7-獆����fn���^Ǘv%��3m�ZxX���H�v�����P�k��mc�D�`��q�鋷�m&����=r��p3d��ڱ��Eyi&��N����̎��(�r�v+���c�}[hm��\n�^�f<�f�HXY=�5�R��FG|B(��%l>��}d2�ۇos�˅}�^�% n��e�m�(��`�-Xc���djh���Sr��SE��ڞ-�B�o�2��@�������[nO. �d�X���"=4�`�
)���)����@��:���9��4W:�]O{��Qa�F���tc������Y���3��Q�>��d_�}�����O��!Q��&�-��+BT�3򒗛��9�	��-�����Z�2�W~���A$��k�a[�9|W�N�&����q����{��H�j�ީ���R�[��D������d|>�dnvnw=�믚*�g���OZ���o����F��;�8��+kµ��$^b�pu3�3���Y5;�Frߘ������t���k>�CMBw�,���F@�ݙ��J�k��e�q��a���w��[��%�A��;�/���oT�/�&����l��䊰h˺D-zM��H��V�m���ג�������3׌ah
��1L͒�w�0�՛��^;8Q�����(S��QO�b��p�M�70��Gp"�9:�
l)@����(jj�^�3�*m՗x�/�:�����	��{��\�|0���?�h<�"��'�sx���J[Q[\���8�w��s�o�wg�ĤvS@\�@��a�[�N�3fcd����>���z8�⾱�摥��7�YWz����.|��ۋ�~���m�և�k?�Sj��ȭ+����{����͓,^��k�:_��U��)_������1�M
��(
�@��7dV:֟ڙ�ax�2�;%|�O��]�%��'?�+m~�`��2Ւx�<����߾�!���m�����u'���gB�%��52��;/�Ag��o�$AuA lTQH��.����/g����~�
z�d����M�j���.I�k����K�
%����ߵU���Í�"�QL0����7VN�����Y4[��۲K�uP��TQ�/�6�-{�h��B�Y�j�_���
nP>�c���3'��A�2��)�a�$��JsJ�-*&���|g��n-�Dc'S�~G	�3��I��T�ڐ�,$���0m�)|�����'W@&�I��X�l���O�6�7F;�*�C���+�W4S!U�Ia�iH.�>1���~]ᨓP֤z$��0"��Jӡ*���l�Q��&K���b��K���Ĵ�U�\� �s��Z=j�P"/���ߕ����^�41c���h�<�*fKH�R��2�¬0���|��p�oGG88*��Ե/�����wP�n6�~|n��lG�9�P���~�BB�3j����z��T��m�����~��\���N���r����Ɖߣ�A���8��ӖэYES'd��R�7@���^�4#b�E��1.�/J$�M����:�[Ng,>i���hTU���N4e8�]���ƞ�_�Og��x=U��k�N��(��_��Ml���hw�"-L�3C�܆�w8f����:$������K(��<�MI�i���ZJ����o�=��0�=��df��^GUNnb"�0i�@��d^�]l�}	+��������!_��7}A3��?�q|�Vo9}�B���.�}Z�L���H��
�1گ�}�tᐝ=��OQ뽃W�����T�@���c������e��t��h}�ODˬ�P�������	d:��w)=�!TwE1�'Nd�9��W��&�i1	�j�;M�2�2I��s��� 2U&n��:���[a����<�k~$�g[oR-��8�ݩ=�6>�\ұmAa�/�1��UF�y�C�`���W�g�"��K��Rj�E�S�~��*3Z���+|��PQ:��'^:����{U�ٿ."0�qb�۰���#�#��1��V(�fB�H�����֬�S�Bۜ$MS4D�@`V�ܬ."��L�VH�? �#�/M때���M	+���%-̱`ͽ�1�Af��!B�{ qH�rP�=+�g8�@8�,(�J��Q��^��N;6���xC�x ��
�+��ϯ(�])�O����U���_aۏY�K"A�P#B�%?��ը]��?��Y���On��IЎu��V!zi���=�*�<���u��p@�ı	-ʄ�e1'��C@����ó����f7���}KȬ�>����k߭j��>`�֧��=|��O�5༌V��؎@˓#[˔p�0�h�S{t'qv�=[���c��a~p�]�ǨS����'pVt_��BF�\����;��ß��(U��LB�#��#�1���.x��v�~xS�N�)" 	;�YEM��U2���?��B(Y`!*�8b'��uz�j��uߴ8�R�-M�I�AOVh3��i���#�*���1�5&1[{GN	��A�gc����%hRT��^B���}j�>�A��-=2fc��ɈJsc�3�.?@]����Е�p�pzt��(��B�i�D�h��4;HB�QFc~�y�)P& �`L�b���i���3�G��\.�iM�sn&��$G���OaX�!��%� ~S���y��ɖu���+g�<(d�$05��(��X�f:�6��A:E�ɷ�+M��2\Ի23[0�F��q��b����7_Ti�j��K����9�W�E~��3wmd	����gޢ�Ʃ�,����	����4)�1n�BN0IM��8;�<�s�p�������UI�1��$(G�U�b�V�^9�O�if{��R��*��yO�0��T&*��+�I�K,	.]|?�ˎ�� t�[���V��9	�\��
��T<�����4
��뺟~<�
Pa��.�D�&I��:��S��p�
�%f�B�*�D��ā��e��""$�|��>�L<E�r�+�X9������'�NqGx��5���x'SR��+��i�2������'g�FV�}u�*�UAۡ�)́�-�x�$�Og�I�����p�V}��}��#��8|�q�OL�~|#���d:i�A����+0��$O���j&��w1��>�Љ��ϳ��?��+����p��¦���?�2ɠ�id��-���;�K��oa@b�K/�>3��=��n[K.�phQ1�?��O'����f������k$��p� P�����t�w��L�7��&&��ђ�(�k�}*�h	��Kˉ�q�'auq����4�����D)��j0�,��iu�v�p`�]	��ڻ�M��Ov�B�iEr�C�U.<�~��JL�3U��l)��'�`(�W-�G,�Xˡ�4��+�;��S<Ғ��������/`<ќ����$�	�� �@vR����+y�=2�:1,���(�/��K�Ӽ�*��،fN�X�ډ�DmDu�(�F����z�
���B�	vw�ڦ�@KO�B���3k����l-f.FX�	JČ�H̀&��f[����?�7���y��.[�{�M�;͚���!�-��2(�J�$�� ز�NSju���Ë���
����޺�R>���¶[��S���0�Q U��������k<��Vn�3b9D�_����LdO>���'+�XCu#�DN��'e�"^���ĲF�A�qG�������Z��4�*&
�ك����6�o��H�%��=}�l,ۈ���{�]���4����i�w������ķξ�Wx�SO��[n��M�U]�.eg��yo(�ZOQ�z���Z��<�x��� ���3EŖ�'�XRH�R�{�x����~�5v'��_��V緔�i�u~|
)�(�lG��^�mZ�U�><2��w
R������?���I'�������+nF�����T��rʄ`-Z1+M��H,��� A8��7
�Sc��,��-���1Z��bh9�[ۘ@����Z��G ���$7<z���Z���/R"/Oޯ"Ę,2��U�k�7Xv}ś�m~�H�OH�i0�!�o���F�Q�VSw�n�*�qp�3�[�����2J?qH~�b���	�Yi\QL��U6)�ŜoɊn4�N�
��u�I���+�$�/D7�b+s*�O-5�fiDm9ū��-ce��;���ll-�_���l���?[��W�Z�+j��
=P���W3ڻN'`I��4�z������=L�?ͽZ�#��6گD��N�sS�/�8ͺ|��<�B��uZy���]�ϋO�����8~�8;�ie�����9q@���jBڀ�K|i$�4���#<�5�:EikQxYp���G�
Ζ�%�)�$���0LǠ�lĕ�����ǓqPE2��A��9����qc���cq�׻��k����;�ԩ�!�xFߍQ5�N��)�GZs�qN�=΄:�Eݲ��������9KT��0�T��[�����q����y<�s4e{ ����BC���y���)��暬���ᐙ���i�D�*���\�.T�n��=��~��?�N��󠌤A��2�ʈM5��Mh5�sy��߷����y��FO����9�I��sk��t��8PZ-��P�~�]A�O�֔�c*����R�P�J6���-"Af��kyQ\�PRXt~�w���y����J#����i'��� ky�e�|B>�sKHR������KH)~�ۙ%9�=�e�Gy�%�9�L�M9��W��+��5�8���C+�k�f��/P��@���H�p���������[c��[4���&�RA6_}�Cda���	�O�|N�g��)u	�n�������xh9�58EzB��˚�j�J��V)z�*��F�o9�E�������.�	,E/C,խC�W���o�mR`3L�*��%��>&��?�0�2BFڊ�㡏����
{��!Ő�^o&P���W!�+<�6t�_כ�����q��G���p>�C���b*AFt�\��ٌ'����lݓ��.W]����u�'�>���z� �3cB��iH�+�J��7�qͺOڜ�ڜB���7�,�qYȟ��M��=�1�%pF ��������ϭ�s9g����ԓP��h������l�]v, Dbe��"@����G�}�^&'/��e���e#�+&!o�帬�@f-Ǔ�
�[@w��a����)��btq�j�&"X?�vzr��n�+/N	��Pq�|sU0�⨌����	��ۡ�)�+T'������.��f>9,=O��',Pq�0ެ=�>itmT�2���LSӽ����z#���]��BXN:�k��n*�0��#F�Z�Ѐ,����7 �g�Ǜ��/Y[��g���EgO��"0�,��_.���=����e��I^��iG�d�����G���rCr����Q��4�M�*fdT�a�O�*]Fؐ�L�E�cmJ?(MN�x{+�g@g�o����W��%.I������oٟ�?Z�j�I���ڴ��e�q'�*^��1�������j�`S��=�q҄)�@5)��~E#����!��EN��6�6�~�!	�������_7!!<v|rk��IG|u �s�ً�gQ�UaX�G�Ӎ�3 �z�6:_���U3��l���y�zD�����zOK+�F��h�%���ݼ��׹;c"���;����ǵ�'7PD�w'�{=��ѓe�x�4}]�&z��Ci� �[���ȕ}�iR���eU:���ԯ�ʹw�%s}%А��.�/F����8�K(À�� 8Ӛ�1VF)��DT��Y[Jp4��WE��O�A�O�&b$o��cJ�v��`�K���Us �j8�߅G:�����Dl�2�hc�� �����׉*֧��O2��;nU_�5BZbFb����EPԗ�ZM��*!�����G]~��"!�	��A9�F�����`��.��nd�����i�t��·�o;JC�f�j��#�_�\mT�Dg-��ʗ.xg�,�W.^����R��h ����qa����˚ֺ��6gn���z�?`'ȍ�j�N�y���`�7D���毱�G��_�69l���Y�~���t@���f��׻�2΍�a_V}	[;�z}|�ֺF��$g��l����f�Q�Iy�r�`�	������PQ���Qar\a�l9�� r\o�̆o��D�C��̛�>� �,_�t
�J��gF�IyE.�g�������℞���k�Հ�z�%�IF��w��F�%��Q.r�S�A�Nz�,��K]Mp	�8��*�gn�?�Ǒ�}<-|�Ǚ��)����cNN�ۼYu�	\�^:&�E)��~T3W��%��c����q��>ђ��Xz����a(���[����jE��{?ҖK:ŕ���)[N�M-O�򳞺;��{��k�EgB�q���w��~%��q�����FE�R�V7Bބ��Q�����)���̬*�BI٫BI�}�w���@��І�Ҫ02�����b<2m;���q������g��%i�����	��?�e��Pғ�zo���ret��n��q�ζr�Vj<��xD�����"�QG;93p���}U4i;�7e����5�ھ-ؤz�k�)^c9�,��h���+S4��N�%"F��l�AD}��N������?eZ�33�K<\��R�]<�<n�hB�3�,���[]��]���|��* =� ��#@��%���J��.�W232���R}m!�)?l���j!U�$��������	+^$��fV�0l�͙@Z�����[ir�@�He3��ҷ�&CDgx�0��<$��(��z���ڰ,rj��?���=dO���{����㉰7��L1�I����O��]����D��< �X<ք�_5/;|n��m{ 7R�Ї9YS����<9L��M�Y)�l�qU-����I�<$U��$��(���#!��ȡ�#&Т���L�U)*��Gˣ#�e�4�	1���`�e8����H�_l���K���d^��'.�i�`��cr�X9�z}S~=,9K�'!���Q�v���~�+_�����h8~��p�W��o�@ț�A��'?]��,~YI�'B�~����S��hOݵ�/c2���KowCϷ�`��:�؁�R���Kj���Gr��/V353,�z>/�!4u�)T-(��O��c�2Hy!H�	"/�5��@�~?U#�4�+8K.7���V����^ٛ*�j)�v������b>2X[J\�P�R��6�C�����B�"H����
.�����:6(�%�� �w�k� ��%�S�ǖC<�V*�\e�(��o+��_Bh-��;���.�3[�w������:�������;�ϳ��+Ҟ�V3���Ϸf�Ϸ�����k;��Y��ŭy�}Ѱ�Z�!2�"�SQ�����Ev��{��)�(�F��9� ��W?yg�[����d�>( ���{d�`��w,�p`�M�rs_z;.:�.���E3�t%B�H840�F�ha��+��?L̝R$=����Iqsω�&CG��g\�su�?u�(��V�3.Z�1���D����=�������W����s��l��q;Fv�Lq�̲e�}ێ��8��JF4l!�!�Ȗ���������u�\.�s����~����u��7�����o��@Ϧ�����%@7��fv)%���s_�p�l�����d'�$H¼�FR�(�9õc�|�bS����1!����@5�x4�&l;�l!���8:��*�:����V]���[U����Z��e3��ϝ�gWh�oK�E�7n�ʘ��Um~:�y�p����9�,lN
|m �vl�z]���0ժc�������x����B́|&�eUQ��1ߙgwsn/3����fm�*���p�he'��;�6��^k�?�'��J�3Q�&E�ll��T���$�,Bx�Ѭ��(.��K��t:8֡r��P}�$#Uā�AH]��S�"��3�!]d���܌��<��~ziBt�4�j�����:r���Y�r2��������h��zѐ�����Ƒ�=!�y��z��HS�b�B���b֓���G��1�h������&���֭��J^7&Å\��"�h��M3ߚ}=���Yя�.�	R��bU�;a9�s>9;�Ӷa�����{�)-��zٕ���Nu�:)f~���'J
>G�6a;�!s4���!��o�w�'x��B��4�c=zuv�NLlY#��Z�2RO���S��}XQ������_��8�#k��B����ܐZ�=2K�_n�s�a��pLʒ���1w�)4[������@�������[�Cj�����ch�S[�TOx��Wb�S�-���7'O��oz�c���֠ݭ�܁��X��[�k�C72���S�Ӭ)���ܒ"������O�6���;q<A��>��D��v�<��!�����L?�����8P]���<$�v��1����6k�Iz����"���e��V������������x�����cL��I��mwM'���]����>8���~nY�|�X}.��Č��$c��<��d�ćXvԣ~��]�����DΛ�18i��Y�����ˡ���w쫈�d�7ɽ]Z�^;�ty��Z���ڄH焬�7��e�=�����+3OD��M���"�$y����㏚L�o�*{��1L��<ӓŪ8^p������H7��8]�9HA����(	/{���/�	���� �~0��x�^�ɸ#����ڻ�mS	G��A$o�*�*b�,��:���s�ӟ��Ù~��4�q&�#��g�z��!B=c��a�x*g��ޕ���R%�� :�4wT�Q���{��7�kǮ�#� �
Z�����Y�,�ʞ��RF��������m��uI��'k�ݼ�g8��(���HnM�`��ˏK�Fˎ����,R�Hx�.P�$�g�!܅F��xj0���f�\C.������fh�a;h���i������Օ7Z�Ov��.E��;:Ot���SYIjbb��nGLn�����b�N�@ݢ�b����D���	YB��������b�G���K�t�9!�7�wV@��Ǘ�u�iw;)M�Ew�Jn5tv��|qY:�������G�|��UQ/��� �e2�=��Iz��g���f}"wm�������ښ���l&5tݏ#�G,)�Q�<���eo�A��Q~�e��]��"�K��viq��~�������հ��<���9V�����ݔH��	�[��� ]�tn�J�ƣ�nLqkj��@�OC�>+2�R�p���Mԃey�K��U�;/��s��Yp^CllM{!��ɂ����T��h"ԥ�<��v��|րF����q%-Ԯ��
�����sjcu[!T�����j���:F:�¸vǨ��,�t�.�X&�&����y�p�&�G�G�R���8K�n�x)�ɷ�m]3=�����������������?:��RA'�6�7���?V�:r�X
<��p~ը�Z�-�j����sZ�GN��G�?�<��	r4���P�{w.�{m��M�'NI5��2�~�<-��+��a��)���R�#��O�E�-�I��m'*��2��U��ؓ�e��
G�o��Zlm�#Y2mZ�7���Y�2C������3כ�g���)=s�_qx.�K�������8��Y��0p6����V�rs��kv��{�0^�<�B���ت��թ����Gt�	��0+ߏK�D�)��4�-�~+���d n������Fk;}y)Y�0�@�F�*3��A��N6rCJA�$#�9V�����#�A�.־]\[�����ə�-`��;���H�wj�[S�B�`�h"�:��+qq�f�2j��Ô�t;Z[�^+V�Y}}v�gL��=�z��=,:�T]��)ZB9L �j�$7t��X��,F�:�h�sb̾���3���&��$k�\_�_w(����P�j����p�ޡkD��TV�@�+P~d�%Gb�C�	�?�ޥ�i��S�q|��;���R�P���`2OgO%�9w'F�_W�:~Z�����!�$�fO�u��%����sŦ�,�"܇� ���@~�ke�,��Gy�\��'��^��U>76V�f(��@g�־TWO�6�]��6r�̰����#L$p����9GP�F��k�ASq��`W�Jq)$�y���q�8�|�=�4/W��2��ي����=�����S�#I���K�T�����Їj�)	�=�B�Z��
ъ'�E��T�nK����s5�}Ij�*w�"�'G1TڕF�T_
��2�LStk�Y*�p�m��-_1��W�aYh������{�w�?�eU��'9�,x,z 5�x��g��I�g�j���������g
S$�>h^��m
f���W���V"]�{�|a���f^ڰHS�d?Y����yW�_���>S9�wt%sP4b�8��^f{%����fl��߳�ξh鼥<k�_\�����'���9����r�Q�7�뙰+7�^ݭ����v'�����V����أ~k��^3�����ˉ�G����D���C�K����NnJ����lXy(�^OU��H���U��)��h�	�{������T�%�F��f�g���kے�<E5�r
���v��;�r�E�?HT���X#Y��*�@�����Q�h��r}~~�Abf���M�ͯ4k�~���Z����0H�~� �~��x�:��[����%�zZ��;�1!�W��[��T�`'G:j@����k��L�/��]��a|<�Ks����!���)�CC��[�Z;�C6�q��@R �f\�˦yQ���w�(u�/&sn��Z�,sw�
d��W�q���c D��.!ݒ������g��Ӹ2X�Ц�[T�P�{�7�;	���P�q4�Ër~��Ϧ:7�=Zz��I�l�Nʃ*�m��2�Us	�*�>�O �/*Fa��4���;:_vuhs�w:�|���D�f[ߔ������� �� �%s�T?��6��~n��C|u3(�������d��u߃[vl|0f�� y���Cx>E�vw��Y:89pA��R�X��\���X�ܣ�j{���F�ȳ�q�P�1;�����STݳ�Q���ÅrH�<TM��[^"�2���k4��.����t�]}h�}:tN8���l�ئC�D�
� A�Eq̸�W�\��=_��STDF۸;
"�Rb�� �B�����,����~�y� �[+�����
8�;�˹�Gq8L��
�����߯��y�5V�!?"#5��lՍ�'|}XLQ�0��~�E�i�t�1��v�L4���y_� ��W�5��.�V��}_����LĲ��&f���NR�G\W��Ɇ�A������=�ߢ���?�G*:p��M��n/�d���2�ޭ��ݬ|Gi<��/kqc��y��*sۜlp���H�0"ˠ��;�c�=�[�|ӧť>���!-�wY"��,���R֢ ![��ro4cu��ـ� �'�I
�>������
R�ga6}4w2�{� ���myY]��B�?�g0Лש���m�hF��lHSc4���N�h^��S�d ����'$fMڧda����f
bhF4���h���T�sܲ�@5
��C���fwM}�E%��Mm�'6��G}9zԭ.3��U��Է�o�yn�`���rX9��8F)\�I��~.�`3�H��]J^yc	HsA�é�������CGF��YV]_��w�!Nr2=�Х�yv�^�!�b@� �uU��c�{%��f����B�1�w��rS�M^�A1��-�U҈�i+�o��/�tD6W��I�c?�v�t�̪���l��|����������dZM�3��:�ȥ�X��jɎ���ݏо2A���_!�d����;x%�[����D�P�,\�C�O\q�ó�$�i&01|i�0ҡ��#�P�8�@fA~�+�du���(�;?��>Z႓I�����{-�N�N,��J����
����A�iR�X>�|;|�{���^V�� 2$	����H� ���X*�68AF72�?H8H�T����ɉ��M�M�g��N�s_[D?��Oڨ
�o�a�[�G�]�)�M��Z-��3k��B�r�����9�GCeV�w� ��S+%+1�0�
�N�t�u�5cS�X#�Y��z�`Zיb�-f���v��ns{g�Q�E������^f�]o�%Յ����)�p~!� 祟Zř�G��-��w�L��X/�T��_���r*?�38Xs�|T	y��;���c��x�L�WTj��sC�
�?E@��z����w,N+i��oy~��I�J�����]�`c��w�o��0��R�v�݋��O��0�8�xO�4�����d�����O?>�bhq��o�cYx��Yr?���������}�xͭ^��ѵI�+��=����!��t��N��jkՓ^*]�`x$���ȧ�L����gl�w٭K�_��hm����
�����ə!�Br��豛�����8J����)�&���p��f�pz���<�u�W�ǁ9��LD�b\�y+�t/Д�]P	,���Ǚ�H]4x6(H�%|�ލ�l�|~����D������ڶy�]+�7�r����i�Đ�u���H�$�����^Rx���$[k��;����J�l��n\��s�M^ '\�#T\�#�ޑ�L+���ht���8	���.�#�ǫp�@�#E��UpC|��tC�tHp�g�z�+����m�I�[�*"Jn��Q{|g0���on�ÕT�G�I�Lr�>T���{\�|+jv��[��� ��w�@1o��|Ě/�:wc�%(�Z�l��c������g�DU=�rX�[�dfAa��l�=���P� �,Й�����oC��=E�GcP�+���>p���� ��� zE����c����xv�a���f\�M�r)H�~�Q%���W�fe�_O���T�z���Ѳ�!�MI4P��Ɣ�h�3tH��s�TB�ěCc��̂�P�3��\8�.�������$S5�h��.,ᳯ�?JL����qi����M�/����Ҡ����C��H�]8�$�j���i�̊��ϙq@��,3�|�H�M��_�v�QrEq�kR@�\n���υ����XQ@gZޘ�(��|:��Ae�82�c�s�B��hf�$fee�y<1-o?OK�co�/��ΎbJ�K�B\ߦ�Z�<s-�G\�Ɠ^��b�����c�a��?��kÈ�j*��\����c�q�nu&����.�Xn�G��o�����Ec5E�1-J<�}�Z���U���+�Mu�3�mOP�`D�g[K7�H�r���]%����F��)�������(�$�	��K/`�xPʒ��U��OL� /�9��u��2����{�������:RP��U��R�޶w������*)VPL~��B]�si��/���v&��пs�_(��$}��� 8� ��j�� ��"��U��嗗�� ��p̸�<+��bQ�=���@O4����:���Rt�|W��N��̫��B__�D3��w+
���Q�Ifg�u�ʭ�so�	[î�m���b{,n���-����Y�0cH�xEM4�����R}z7��"�r����z�]�?yT6���5�
��k���;��h��5ݼW	T`;W.��#r��iH��L��_�\?]��o�4#0^��+�Et�	BE�2�t(9�)����է�u��.O��ꔮ�D_��.&�����V�3�D&s.��"$ϔbb��,7=Qqb���I+%�+���e7:!Y���"��VDr}qʥ��E t�������}��|:�E)��p�I8����mܲ�w�_^v��@�]��2���L���(D��Rֵ�ud]ʾ����v�
%�-Z'���:ƫwa�������,l���ƫ\`�g�����RD�r��C�+���}��lJߏ�F���,�kHf Aw�+�T!�a��%�DVt�e�'��S2m
��^�="�4^Mg�B&������%���}�b���ɏ����>o��}V�b�u0�k2��<�좂�b�{?Lr���^V8��:�Ei'��#��*�
����H�����=pn��?zK:Y�F��(�sk�K(�T����3��n���m��r��j�]r�z>�̊~V���]��8|�Y6��&Yx�M,���@�I���t��V��$x�a������D^YW^P�=�!� V�xd�A�f��u/yW���W[��`	��3�9�W��!��t��;���i��Zs�c�+�.jh�#��줁��r}�
>(��y&H1^�PX���i��%/=�D7T\Vؔ���4]2w�6��S� 6�:vPZ���Z�yw�������Jh���S�v��>�����O����I'�B��"pQeW�T-d��GO�c/D@����{p�c~�Y�/����	� �@�k��[E�bi���q��Ŷ���s�b��'
'E.^cQ����k�wD|���d��zMi���F�o��_݅�Q
-��=C�O�n��_ǣ�H{O_{��%IѠ��g�E�5,����Q�ľ�d���ȺW�e.n�8z���Տ����SA���0�t)VZ���@Y�`:[q���������(�/~��{۞��֜��l�.m�ᓧ��ٲ@�4�i��o�??���E_��}�V��g�1�U>=��q��ʅ��U���n�N��|!�Z�4s���v(
�FoX1;�,��E���,�`�[��x����ΞmJ���s|ͷ������@at�%�:���i;�ʨ$�8�t���~E�Jl��X���n��w:��L�	�`
̼�m��@>c���b�+�C��G�d�^²v��������L,o���ç,Y:}آp,��7�@���Lm㞸�^�|�h��RX��aG��ri�_pOP*Vn��~���$�#9ʬp��A�O�b�!>ϸ.���9�o�v���ҍ3��7�?��\$�BX�?\�Sfҩ����"g�*|�|$'D>	� ��$��s>r�K-�7x�0�1T�oj�OZ�V���.v����,Uh�������A��}�}���B�ZH���k2�絬13z�\�V�тg~E.7���.��>/ ?�Z����\\~S��ν�<� ���œ�,�K���jƲ�kR��2�0���>:ҥ��x����o�2C䛗��-� [�q"R��uh�sA���Ǆ�P^h�Nm库&[��M8���~�rUS[X)c(Jɐ�����s!�ql�����J�f�a�oǧ�w�(�<���rW�L�OW��P/
�gy��c������I��ϭ����tʍt
�.����-P~�4�����l�� ���Vis��h����%��𥙲���P�o\�5��${����f��������zx]��?A�浕K�֢�`�W�k�/d��̆����N�/�3�\{�Y����И��oi�N��H5��Тb�]���U�b;��^�����0"jj���K��D�t&Ww�tj�tdNL�'B]�<���!��ڜ��,~��58�i{i�ㅻC9�^�F_�.Р�0+~;���,�B@����	e*�y�<�_���z~���B�-���'&�YP�a[�t�W���K<M�8TR�*
�y�ok��슌��3垖y8���=+�<,�����:܅uT��m�'��X
� ���'Ѳ��Ι�m�7�����?r��
�����4<o�ok���<��;^��@y0�_�2$�3\��(���*�ZR�(�=��9���Z�Rv%z�~^�������5C��&����$���7�Hwp�Z�+��\*K��K|T���k\܍��v1�1�c�>�0ղ�7_ N�^+:c�WK�)�˿g��Qw
��yL|f�^ϵ��>�w:�Ӆ�0M��x=6�Ad�)��ma���wF+���q��%g�/��>~�ݩ�<�=��1�)�i��2$�x�ͱ��6��-,z!�K/�u�)ݭK��!�|2#]�#�H��d�Otos��#}��7���zg�NVz���J����X1wrk���u
�����q���K�����*)\7���[j]�.3IM�!�Ab�&!��x����"���d����:}c�߲�^|���B�vn��q
؞K�E3�� ��[-���u��i��[Dx�9V����,25�� 6"�<�RH����vƈ^A��qC+|@]=@Z�h�<.}��:x��0�4��ǆ���O��p��z�$tƥHo7��	��z���)�S�~RZ#O:��w�{�6d����s��~���6���(����$�XC�[['w�� ����.���.�������(�ټ�H��\�\�n�c<5���3�8�80 ma��V���,3@�l�FH�U��*�\��5��L-�a��_��hv�8}Uf�-×�[,_¸�k�-o�>��ge�O�ʨ��/P��[�"�?��J�g �Y�}�;l��$�Dzr�Q�B�8;�/ AFf*��+l0[\�M���.��z��29e��#S3�ә&�����	CDY�R�����n���_bg{0d�s癩���k�=���6K�O���O�v�S��`>�=�el�b1���� ��8{�?���P�r���X7��͐��W�~��z�8����H�o�8R[#��VT���"#IO]�V'��X�dg'���dޕ�[����jp�^�"�i�li��\_i(�����~�#VB� M@fq��58늸C/�n|U�~^J� ˑT,f$�iZ�"�B��]߁����H�z�Q��M���8�lk����V��%E��V�%���gY�g �?,K
h۵�8��^����ˁ�,F��>|��N��A�;�@��4����9=�Jw���͸cEϊ\�DV?#C��5^����:���y�V��F����e���Ʋ����%p��"[��
 ��PĲˋ�O�:��X���N[��UOa�#\��v=yތ�k������=,��֥�.��/�c��������+��]�bs�X�xx��'�r��lj�̡s����`�\r�����O0W�	��pV�v��b�]��������R�l�n��2x����O��k�o@���q�g����U��n�;OI��~�c���Ʉ�p'JDkp�v�ձ^k�ZV��,�AZ(�����bE˺&�Y.� ��J�j�bυ�T��*~}�"ŴW��^��&�&��rTf��dC��x�ǥfE�<G����)�S.�l��^�B.�we�S���~5��k߼�Ռ�

m,�m�s|?Z��FQ��e�)�����d8��h�K�>z��/`�S*�<��a>�f;��ޣ3U�y��ǅDC?:�5cT��O�h"�3�t��(5��)���$;�ВIU@wɥpmy��m|?=��׊ڵ(��=��bp"�(�d }��` -�^��&��҄��_^9��ÈpU�Y���~�����M��.��Y����g��|��.㝧.`�ѐc�~��z�!������D�/~z��qSH,��yq�d�
�F���ݏ;x%�Ry�?p��y	~%���ܾ��	��93�&�;��h!�����3�k�6�S�&��a������HՍ�ЕOw�g��4^�XPC瘑~%VRfnF�3ַ���@� �Ҫ�6e��)܅F����NW�I{Q%�n�p�0?-^��pI�v�v�J���%�L��Uy`Y�")�u�W�,�gk��[`&�iPZL�E����+�Y0�h�Q�a�.���a���pe���˾X��B�̥1/�'�w B Ζ_s�1��G�9i��W<^B�&�	������t���,�l�11�Ѡm��oX��h��b�H|���n��0�$����{z(8�*h<W�Pb|��~�3`�\G%O��L�!��Zõ�k��T��E�ϵ��&hH0���v��|������Eˍ����#�F�6��|��].����S�O3-MW�\�c~�|�DO�מ�4(�"`�HҠ��f���JƱ�T��P�4�2�SJ>�$�
��ERZ����e-ԁ2���d9�����S�&�F�I%/�9Jg8�%�h�H��83��N���b]�������������0FqFJ~>󵉗���,�q`�jD���*�'�>�E�;��NnsJ�����&��7�tdX
/R�2mv҄:�wI��q�%���e+4@�����g��7�w������*�4]'Ov��$�<�
�((հ�'$��c�!<�di��G��������.����D�S3r���m���۱E)�8�����Кh�{"��y��quh����Gq���}�r�*�L2=;���@$�-� ����aK�(�� i���.������H+!u�����J�6W uk����]j��rM<޿�{���Ɨ�sMhB/w��"GO���lj�*n�'+����2��O�zh]a������.Kqތ5�̊pu�D£��b����*�{{:2��K������b��'�{\q��󒪹��h�4��������q����dEc翅)�A"��ņ�[��J��
�L��3���$���u����M=�9��/D�w9�����^'U����ō���t�ĳ�&�f��j:#�g|�M�y	=8���m�8L�ʽa�=F�����+��W\[h݌>%lw(��[���Y�̝�{i�+r�80�-�@�T�'�h����h,��A��S ���E6�9�i�g�^��»Z֓�ޣ�p$�o�?���g�q��.��n���SrqK�H�HC[���Q�[����PiDP�^#�P%V���Ś'H��%ҵ��gB�Ω�_�,#O�P���:I��i 8=�L	F$����2W{vz�����;�Ӿ�f�ϭ����"�U������G���F�K
����|�� v�y�|�az�����,HҐ��d�1s��D��Qմ"���@�Rm�n����'�-C��c)��Ϳ-P�Qd���9�BA����#YL>��Fm�sN��\��%�܏��z�7��	��N���G[�������"��*���Z+�d I1�~��Ԩ�Ood&ɲ����s+�XŦH˙n�(�
'���r�S����@�ݒDϬ��i��>���Ж��'�Pq)���?�
���Fm�>ғc@:�h�xh��T]�L�����{���l6CsH�#����'��,�]�w�;Q�h�'�!��Y�z��ha���cWE�.�E���1Gl�R�$VF�*���Y��q�����(�v%Z��0hUR�r4a��ԕ(��n*s	ʡ�D�\R��~���ӋE��fTY�V��˦��~�AN��^<�����fp�����f�<��f̀��侰�[�:��!U�v^b?�	���N��?����u�'��,���%�Ǚ�j@�����Pi�0;���M�NKĩ��`��=��
�(�*E��<� �$�ЮJ�,
����m�
�ݫ�T�\����)�����, ~'Y0*���+?8%�YAA�=$����ê�ܪ[E:
͔�6���ZWajHISbû��go�+�\�*�
c^���N�"����Olw�q��x홉����U�gR��4$�����8: �<���֪��<�F��C�5.��^W5�%�f�$<�u�YYVU�k�?W�CC|w��[U���5�Z����Q%��뒅��T_'ޱ�I6/I�ل���,$�os�6r���zz)��.S(�to6��[<+�3�1��k͇c����}n�k�FD&��A��ﾫ�l*8�|�-��A��x��58�5��7k�(6^����u�[��~�w?�da�,U���#ƀf,��w�s� �%�+�x��2.��`��EHv��� -;`�/���Mԃ��}(�%Qbg5�P=B u��b��[��T�M7\a��%��c��/��5-h��+4SN��mU�ig�ߟ�Y����Z�3E
E��zp��MԋP[��/�t1��.E��x�j�ց.ŋ���B@T��ֺC}�nJT���\����'v��$�G�Ňto�uz��;(�U�.�2��\Hum��=�8��o�a]����}9�D��B�>�WO	����"�(z��,��R������6����f����*�v�9P��3`����pԬ����޺�ˊ��d���eZ���ܝ���������w�����t`G98�w�* ă'm-s�h�Fda��؉JV:���bz"���e�HkԷo*�`�|+5�B�j6��Bq�;9�ҹS�ٟ�~*�O;t7��3\�s䅜.��׼�������ǥ�|ѥ�ᚙ��&��.���+$%�q�_�@��>����$���/Zlb�֓hF��Is ك��K�� 7�&r`k�����3���8������֩�x��f��{�:�8ϼDn���E��<����ւ(4�5�OR�	�~H��!]�����=bE �҇b&�W����G�x2�����S��Kx46M��`e�؅��%��i��?sX�%p���nQq7$.HQ����F�O�60'�k^�� V\&��f�q����%�a����pA.R>6	��)�so΃KU7���yUpi��ب:/��yp,C���w�'41�e�D3��P0�i:�	\�
i*吭8�@�7���duO��Tyu�E$�)�����۟���a�h@��wae
a��C.����:6�ᐡ�W�Y�QA���陴&$�_�����ΰ�0J�!zc3JW+��Q�#�7޿q�M���!����/�����S�"3Xa˿�58�.�_oIC$��d�xd� {j8�\��6Ġ*ާ����j4�L�~	��1��:�\�'���$Mm�ɮ��gﭑ�S�4=	P���;d�pr�Y�k ��7o3�rP�fN���JJy	^-���8��Z�>/8�m@k��E?��癖��c�%���g'#��6�������� �����:J?J[��?���~C{�Һ�&��0���W����
�a��S�]P�9�I]���%����"��U<{���
,�8c�|o�W`��Ul�3�-����p-6��{	�X�66M���|���	G6A�l��iz�<iک�tD̵隉�l���C��R	�D[+<�c�-.nlr5���i�pa�,(�T���h�j^�Ϲyw7�-gӏN��A��ݻ�[��vs?�ߏ�	0k-nK�����zL	���X�J)��s��jӶ����y�[�=��O5�څ�Ns�o��� H�����)� �d ��H�AaJ�\^�U�UI��X�ӈ���8�e�p9J�_�hR�y@ܑ��m�!;���J�Ub,ah�m�"/r{}�b<q�I\����m���P������5�AC�9�~�_x��]g��m��.�뻋�����=.F�[���X�l�_j��_'���CODZ�zq��y�w��A�"\��P�B�La9D�,���R�_A��LS_!Һ�ϓ���]a��s�2#��e����x��gП��t��IƙΌ�7.��j+��ygݢ6F�L��W����.�hS�%pQobD�}|˟uO������fU�d��g羛R#�_�$�0��� �C��BDr�=�3Su�qmO��5/�� ����ο7��xX����S�%4�rS�Ӟ����ө�H���/n8Fi�5�`"RmzŊP9�Fr���/V��\u�@W=��Z��Wjc�P�7����bλXkB�妀�ף�HCU�����C�'�0ً�;)�}�njƝl��	�tR�d�����P������4�Q�~�Zq�4��8�~�^�t�w���ӌ��كc���O��i�r�����W���	�H88r�#�j�9�����\j`�*�
6Y�姂$'\6�LLlkZ��|�G�J�:҂k� ��Otv��`��ѿ.�M��#6�|'��+�j`��TB|W���uW��W����M�5�^�7�\J���؟p |Ő��Uv��	��P�΃��Θs�j��pr�%�+�-*6k�6`7����:ԟ荭��M/��0���v�R��p��x	�"��E8�d�_�HB
��E	L*�/r�W���N��;������`z?���§�.���ܯb�ڇ{O���]����y+�(�}u����Rh��rG�🌶X"i���F�r
ٲ�R���F�Y��]	xp�c�<��x�t�:�Y�B8uT�+��,�k��*�++��GD����܄x���0�[4��9��u�������Фe&��r	�4�W��$��(�ؗG�L���|�^���W���;��@�5BuJHWaP?�$@�ҭ-r��5ͺX��(�l�.d�b	��Y��E<�j �cWjLszsIaz��qWЏ�Q���
����Wok�,\?�D-���r�^�f��|"� D�{�����F٦��ں���1CH�dC��آwe�H���.A�e�7���gd�6��+^v�pc�zX_)�l�>���IV�(��Zt���Ʌur+a�����l�2��:�m�2�Q�p~&�����t��j�6g=���ה����&��%G*���g���7؄xU�ͱ�SI���X���)㿖�26�?�����ߟV�ګ�3�89~=���No?,������K���{o\����
R})�]��)0)�ɕ��M?�f�N9a�/��+v�Q��E�8��O²�.<�NB�_��тY~2�Ÿ|�i�1��Rr���݆m���0��%���w�&P��@��O��(ǈ�E���|^+a������6Q����uɻJ���!��x�e��'���O}�YJ]�"߄��6,;hn����Y���"�H���v�594>6Y=���7����	���a��N�����!1v�/��>�Y���*=氻�̊�S��A�/�9o~$��./w\s����@Y����ϗ��{ڧ��q:��FK'&jܭ����e�g�H�qO��T렙ō��B{
��&���� ���m��d�� _���>ױW�gL�Q4��o�!1���F���BsC'#�,����F�2C�0�;U����m�;ȕ�g���kBY}X�fa��������0��źLw�
��)�3�q�M-�Gr[��L���4�o+�e%<|�ni\�� ������i�hd��p~�A�k×
PV�I�e���/
��?�M� zb#6��_��2�J��:P�'x�qs�B/�dV�(E�P�+/E��P�N�J��,}���}�T�T��op�X��8g.nCV� �A��נ�b�f�_ 2w����S�3�s���G����͘<V����3��c7U���U֗,c7�\���?���d)X4O�e)�Ì�c(X����w�F�U9M���.zȮ��ϳ��j����'~{��R��ȁ������b�n,)+)"1����W��>I�x�*�fk?����geG��|FQ������b$�+�B��@�oJ�Q������%:\/�T-}��2�ӑ�?ɉT��M �	g��ꎷ}�cg������*ѳQ�.���R�Ե/�w�����G�Lm,$�f�}d�T�"���W"�I-��b�l�o�i^���~UbkZUq��
sNn�͡Q&p%e[�s:���IZɋSŧ]B- ):b�;z��1��q-�&��ԟ�Š�����J-����Fw}����biI��J��G���Ql�GT�� O��h�)��
�c���ߌ�fK���S�Y�	L�(����a˩����\� �s+\�FJ��b�*D���h�a��gv�OK���y��P�CU0ɵ�&�Iok(&yD�c�?�y��?�cr7=jiݚ�&A>W'-��d�b�N����碲�_�N���t�����A�i��^��_�D1yV�#�Rܯ��VV�Y����^R��(>V��J9��I�H����r/צ��U�!���1^����H�!M��\u���%/�5��sEA)xϞ�H� R����î�5f�+�7�yX]&�,�4���c�OY�"��6���{xT�d�5_����s��l,}�e�w����y1ցw]T�S���
���;Q	D<r�Gw7Ǌ��R	2況,]�p�S�m�Y\�E����">�OWԵ����w/ސ��X${֊Ѵ��
H��B�g�w�۞��δ�?},�#�9��p��1����]������NDF5Z��.�0�'����Q}fb�\�Q��R��9 �hpm{\���"̀6׼��yb��!���#��t~kPl�9���"6}�DX��� ���7�@��?��1z³��o�~:oӊ�z~������aM�a��R���0��0F�0JPB:D���p�hF7:DRR�*�-�H# -!���>��}��yw��{��s�y��u���;;��52�����B]��O��:��|S�]��/ 2ம.ε�������c�fq��2��}b�ۜ[�IUN�M[�����5ʽ���{�q���$`�K�'+5"ϵ����Ђ��7���.'�`���(����S>q�w���'}��ާ#�d�%�~�V�l��:��
^JeT�Z�z�~t�
��Sy��o�p�'r�E��N�E��A���N~r�����/3�弛%���	)�K!L���W�����
����-��A٭�X0|�N����p�a�2=��9�zx�f�Ɏ+115� ������u��oVb�~��&��"Iٿ6N�[���n���2Ό�o�h��3�Q!�������&��q�5�`w�oqT�Ĕ~��H͐d9�Rw�=w�)��)�R|܈�AS�2�VHԉNW~�b��}B�����{����=����"��EulDq<�Kn���H�5����P}������2Xm�?��J��j��Q��[(&�C_녳�M�#��fx�B���[%R~���kq����cߔ�ED�)}}>��+��V`_ �tK� �n~"�����E��a��OmVH3/Ƽ�I�k���=G��*���F����*�ۮ�%+`����^O��?����@Ub�}����L5LUGMK��.#UJ5�}_�b�HhH d��y� �n	��P�
"1�]��1�ox|_�sj��+;�(�~�m[��fᔉ�(<5 6�"��?��{�2kӞvG�
�w���@�ze�)L����C��8��G&Mۚ�@1�m"q:0�g�v�@���"q*I���)HLǄ��>����Y@�=Z!��PsӜ)��������l����9��S�4�By)R��q���W���S�ܯ|�`��W+���t����KZ�I��&rG��B9�������X�<��r���(��Nk�����g@�Ӈ��\�a���0I���޷�U1ĥ��x�9ɘ��?�^"e6�ىuT2'y*��^�ǝ'w�+�4b}Cm3.�^�d�j�0�&eJ�:h��O��Ԡ�Aن���������-�i=Ht%hL@�F/�W�;�A�Ԕ�³� 6Z��雮��������$l�l=�=!ؚ�1� ]�ޒ4A�b�k`�.�D�b�r�v�����
��M3��0�@�[j�{����OO��!֩Wl(���XB�Z�t�:h��jc�u��ͮ��Zt������Y�CX�t:3`�#!���;TDb�S&/��Z�.`�_�Z5XX4n��u���wL.󭞶]��fS��P�[^9�С2�_D,T���KͿh�oz��}<��� 6~����K		o�o���Z��P`�����u�q0	6+$�O�f��(^�DX=b�J��_	H?;o�殥���<dS8�+�C��b{H{h��زz>����y^�� ����"t���z�۸���J�d��3�Rjߞ���z�,1z��g�����H`O��"V������gw.�ׅ��L�x�=��K+�#��B ٛ0�P�}���b�Əb����!���ٷ�B��p{�-@��d�3#�B�^GE��U��u=�)��f/���p�9�60���˖�T�n+"�P���fa	��q�g-ɛ��FC
�ݷj�5 _�4	r�>R�nC����n{�:�
��y��?��A�ej�N����H/��PO#��������I-�/0h��~jGL�'����5U���r����ol�U}�Gє�3ȓ-�Z>ݢ9�*�Ou�?'R�=o�7006$d$��bp��r��Eʲ�sܜRiF�%@�0�}>�n�	4+Xh7��x��W��M֦�_�vK'����{:<q��^'Z��W�\7x�5O��xA1��$��ig�>\����Mݕ���5�o�����M��Fy&��K)4���j�?�\�pc�5���I�fD�vש��x.����@0����:?:�����i���ր<"0P>�=7]o�p�ޚ�d�\��QI�5�����}�.g�y�A3<>f�_�,��	P���x2��5hk�.L�0��K�Oe�xT���~o[\��M����p�Ge*�zhy?W3{q�{/��n�B��ɫ����i�a$X�u��X��S�N�"��I��W�)��
wƚBR�i*���d��]����/_�\S >��'o��{2�|,�+����#�`�;���2��S��0�����&� �d��B��7�IM�P*�jfI0��Tj[2	�"t���)L���dUC�~;OG�`@�si|��Bb*k>�Xd.��<������;�_e�΂V�Y�R�wM���DHY���G�>�m#N�4]1Q�\3cLj�,5�E�뉚���nE�R��4�T���j8���^�f#��~�{\$Сz:�#���mA����D8�=Ƭ��E5^}2�j��G�N��Z����.��aJ-(o9C��,����<%:���-�
�lkG�>M	"�3b����k���@�p��ߜ��bC:����ĕ
�ɏ����5���]���'up6秦��>���~&�h��{�P�؅H����J��<U&{�y�nX���C��k2���P�T�T
Lǭ\b��.�H��
�p�Y y\Cn}e� �S�Foq����3�P�0�5~`$/Y�~Eo�%���@��f��;]+
�~3p�³?�:{6w��z��]t�ઊ�]�_�v.EB�_��Mh�t��n�-U ,l#�菷{<��(��-{���bù�}�����&���]��8�u2&����EM��5�����ܼ�GW�����A��RԜ�EhgggO��Ĕw�F�^��84���	�^=67�*��L.]����c�� �:H-�D3����ǔ����k�Gw�{:;�Y�F����w�%Ć`(��^r��g�Yu!��>�R�i�|+7�����l��O��dY٠�On�_X}��'��w{7��\�z0 ���9�4r�,�	p��kT-�dBx��oL�Gtƕ�7��$B��ٚ3�W>�2��ӓ,��H�a*��U9�~{��aﭔ�A�^���L�Y����OӲ>j�$ItÎ��K4�L�RdIj/O���h�����bhu9����D�l	nݡ�8���^�}w�[w�;���U�(�EJ�(r>-q�yf�hG)�`s!��K���{mmk40���Hy�������HՐ'�.��8���=3cD\�h4
2�����c�mĸL���Iʡٌ����9�+=�����.�w�,���%f{�wI(Zv��pSRwQ��Q��)�i��C->���CΉH��n����@5N����n��2�c�|�4�)v��ռUixh��9�g��N�ӽm��9t�����^B�Z�t�hTO�{@����v�0���?
!v������>�Vt�f�g{(�X�7Phcq���}#����:�K��ԕ֣��[��p}ypH=y�W�KfA=�ɥC���+<
l�"�B��L��A��@RD����n�ؤ+٧߭!��ru�W�&�uV�*�5"v4"��!iqZk���qL{���>.&0��Z��*�T=�ud������!�p��~�9}lS����0ǹJ�wo^��-�}Po~���4`����ޮ	B�-j�/'�{����,O��> ,h��D�m@�ʊ>Ӥ�tP�F���L�,��I�����IKǕ��.,��N�NE��r��_
#K-��c�A��������.?2w~���Z�vE�p�oo����u�+�������ǁL�:��f�g��A�&��uaF��*^���*Z��īEs���"�P�_�m n��h���萞���F

�4K_�
�pz���24Z��^�u�X\K�G��@mg����'Faj鸐����Q�~�WK�Q�bJ�����-��>�ݽ��Tzi�'�i�yɯ�a��3�P����q�d��1 +���w����w��jb�� �$U���y� ���asqz�R��K5��»"Ѱ��gp��+��L��n��=�mK���E8�����;T8���*��NU���BЃ�R��Q��I�X�@��_�G>�܄���G	�L=[�y_��	�_{���8���+j9�g?;C��&̜+1�;�Y��.1�sQ%�'
ه�3��y�Jů��2�2�{!\��(V� �8�������~?��MG ���e�g&;��׵W�el(�5�&l�Q'˺uGO�-��0��v�'(�N�7��=�k�z�TC���Y�ed������P'ŷC�T�.t@L�ӣ,[JK@ ��[���LI+�wi�����w�/HP���/v,'?�����A j�%�WD5}�.6� �
�Q�����	O��L:w��Y�A��2�j'��m>l~�{���L�	Q�:x�?����"�ON���QFĔQ��6�OOtuz���+0��|A�a�:�ȝ�' FF��q������s��/��/�<�
���~���U���E��f�-a�s�bk�d����=Q��U@���� j# j&@��c�}LY����ƷqАR����P.`�(����^�N�_��"��$Ѩ�P���2O\�1&z�nJ8�+�T��!l�	�hȏ�S�����ǵ98�
�8�����-����F�J]x����/�^�h/"���ewl��##)6&�kb8��1<���̓	�,q=�֩x�@ZR��e"u�٣�?�<�E�z���!Pd\�ZI�:��~9ۢ�
�8-���IK�G�E�|�fsl�}b�T�0��A�l���i9h?���"qN�qn���]p�oᤤ.zo3ƶ�4`'5$ݲ��k���M����W�Ĉ�r���绐�h��{�PB�*��Ҁ�0���<�m;�
�(T�|��']�@_�kŶ,��FY򲡺���K��?�8���R�P�������;$���g��5I[Z�
f�?/Y�=�\�]��[�Ν>�Ч��Ճ������������Yե��?�4{��⣇Q$�	� �EhØJ1�B˔
!������$�P��us^�/��@�� +&��g(�E$=Ø@3?aY+�9���{�~kU���H��R��Wߥ{g�7o�Ѣ3�����mu�K��bd����{꼩�����O�M����p?*���b�P�'�3 �g���I��9TU��K�gn}�)�+������%����[!��탥���#΀|���	ib�]��7��|&�>n9�V���I�����CL^.�z"�
�����߼�"7�aʗ��`�k�n��D�e�u�X�)1l	�J*���bi�+�=Y7
�z*�����yJζl�Igp�{��$��m{����.��<.
��^*��:�`'	Iv�8I`��|���V,��wN���o٨�Kh\	Uq����&����1��:�MMaH�"ޘD�ups���$�T��-꤭�T�Zz�؆{��0�":/�9�Ϸ��- �;6:I����ol�bp�V����'��~��腙Of�{��M
2>�&��I�z2_�׶Z�-� ���:A����28ݭ�#��Ӯ4V$צO0�We�OJ�bg1�A\�셅_[�F
�u݂|T��bC��9���
�y`��`&T�J~��-v�~��5���j���V�)��Ҁ��Ly�|O�P
U�N�����ϗ���KA�if�:(��b?~ږv�9{Kf�,䐚�i2�E��=�fij�'�t,=#��qA
~RC�D��9q%�^Nw�`,j���3��c�
��(\է2�qblÀꄅ�<�a��i���D(���\��r��ўyv�@1��KA�(T�)T���0D}KF�p@�� �L��������m���e:�1c�ȃ`%��P��g`@�����s�Y��Q���N(�j;C�8݆����;�j��8W}﯀b�6O���4�|GP�F	�*V�J���ox� �K�#F.�C �3��_���y�rl�E�����ģ )�a)�����p{��|5�UjWFf���{yUR=�d�'56���}Ϡ�s���2�����@yGL�{V�O ����r�t��eg9�Q8��O������/!(X�y��2��h�P��2�H� ��*$٫S{$j�����cBE����Z��\�pv[���-.���d�h�=ه?���2ry{��1MvJ�;4B��g�ظ�o���%D !��DL��:����ShR�e��X����H�Qg�Vk'_샎�50:��[No�l�Ƹ�
�'��俉>!!��^�}Ku�����K9�Aq(�B�D��Fy=�F� ���J�e����[�����5�P�"ԉ_j�D;��(]��H��c�vgKbo�\xrW��7�+��V!3��t's��ug ���&�B��kO5I�7��/&�m\N/�}RRFi{���Sxv)_�y#W���k0F��K-3U����3�_A.Ww�X�Z���j)A���&l@L)�pk8ርc'����d+9�-Y�g�TY�9[F17�-7�"�!ވ]�����酹�]osd@ѫ��F��~��Ц~m��x" ,aU� 7�6a�Ҳ0�~%3pB�*��0�>�Y1��-y�lJ�VJ���uP>��*��f��$0tk�r 4x+Ӝ�Fv����,e�we���:�5���!<�+�ݠ��E�_�kn�3��ݔ=�!�����*Q��X^�wu��U~Δ&ͩ��[J�Ve»�4��M����I��'��NO��'',��({v=B�WZ�,��G��+�ٖ*�Л��������ܾ�+W"��	x��{m�I���)CU���3�N�{�*�K��j�I��Z4C9eS:N�I��	�&�E�K�B��dj:Hx��8[%#����Dӟ��k �ѫ����Ex��D��R�{C1�����ql�������=l��1O�Rp���@oo��0E��cf}5Ƞ/�ء��)��1�2�@o�̋�  �Ċ�U(G���	���B2�ٯ4d��3�!u�S�m �����4�yM��Ԙ�j���'k�-��J����yz(��^W��;|�}��� �1�d;���e�Qp��׃���边A��\f�+���@��b�xrf9)��ϴ��J$�>���W��O�Ӏn$F��v�-޿௮��H��/GBc�$r���!Z�@����8�H<��̾v|��]}qw+��V���{����O�^�k��
�[����5����.y���;' ��F<��P���� ��LǄ>*�)�UĐi�)��o�*�X�ﭓL�1JY�m=i,l�,U�=\�)���Q%%�p�O\ܓ�	��ʚ�ً��@��W{�\u��0�՘K��=TBb�:��f��K �N��ҿOr,�T�zbF[t
7���ˡ$��=�-\)Ȧ�#j3��~� 9&�	�uU��S��7��'T��7S�}�&�G�3EmZ������5�u#k����UdԞS�����>�O&ɴ����;���,�}ۈW��~j�L�y��/A��D!���,����������ќ�i�d�L��*5k�9���U��^���v�EZ�,��=�H�=�I���a�6�w�O�O�*���d)^?HN���w��r��q�
�T��J�~������gύT�H��T�W�������-9nF9o����tN��m��������t�V���)�@Mxe��fgÈ�Dq��A@�[5%(�5�m���g�?��ۻ�rGXft�A���$V Κ�P|}�vh����g^�0X�5�u��&��Kz�W�7S��_�*���~����|q�*�C�eO��9���ć�#ۢ��5��S�#�՜��~7|j�Ɏ�K����	���}�?;Z��������C��<����Q�bAr��A���!�b�s���m++6fQۄS�V������Fjn�Q���zg�0�@�L��&mX��P�R�2�
�3�G1��ʳ��[��|O>7�'�P�,P�,��m>�ӫ����;�Zd~�f����x�����!����b�3�b��H@�f(��j�	����Ա+2qƛ����2&B������M;�4Q��!�6��g vq�����xv�7ϣ��9����Z�z�:�ή�U��&��f�`d�%@ؐ�Sg��̔J$>�]�5��?�=�C�-D��Y�/�gÅ]?+X[P�O�'�4�C1��Y)�5����0��Mg�2��omdo��U{���L��-h���1�9��k꿘��b;;��\������t��;-`���ޙ�U�ӛ � U 5H4aF5+�N'}�"�J�>S�J��B֗e�/3�+�@�ah����t�v����w����$K�3�91t.�^2">����t�H��v�H�+����E�������X��,t�����%��N]��td�N	�P~��j�Ј�J밦����u+j�$�|��o��:`|���oE)2.#��^�c��c��ң��߉��J���?�Z:���O-5���^�W�eځ�]-�F�W�=���	�4Y��C���U6����<rJ7;��YoNƎ��.���ڊm9���v�u�vn��Y��t�l���t�n#����|��چ��;,b���]���L����1�.f�Yijj�A@��m�1�a�����<�T(�� I�����0YlP�C�	%ܗ2��DiH<���2�,�P��n_�a�(�9��5��Aa�Vs5Lⓐ�yvd��{2����W���������W�Al�;5�/J��=��Ǐ�&bGN��_�-���4���s<�ɾ��w�!��!�1_�����½��4�>[K�Y��cw3��D�I�Z�V���Pf� �dz��������l��E-ȝ%��|��ۗ"���j	�B�lw+A�9�/��If$�ݑ��$�>�k��;���0�ࣦ���N��� ��M�x��a����y5_%�ZQ������$wɏ��:q�p*��d`�nۮ����UN�m�BH��{�П��R(%� ����H)��އ2ya>0m2hJ��4v��ą:mȨ���Կ�'�̄�L�����VG�����bH�?Lw;��`��{t����ö)e�X�rP�f�7S��� ���oI_�_a?�.��萃C��g9�!a^�O��ش��H�}�E>�8�;�¢WoM����M�շ�ݹm���C�����������75�O-P�PI���u����|�1�?����|�@�w��u�uZ�W%ML99��4�r��Q����>�O�L��n&����Ē��0���՛�U{����"�e� d7����<����y��@R-P&q��a���.p�L���ٺ}��.��<�����N��}�<��V
�� �4���G�砽�E�s�V�y����m�?2��ܢ"G�`;��N�f� y�f�<���9�rg��Wi=5+���}�z�c����(tO���GH	�ڄ�-��|�9.�K���zG��)Yo�y5����|�#:��;�z���Wm�1��:��.��q^E�ah��.Tز�їE�m�`�I�%�I�nҔ���va���9�q�����8���:I�[Ϩ{�~KM0��A�ޒ�V�ZX�Y�=��!�.���)��[����cj�A5��4���Y�>V	v6(BP�
��<h�D���5�v{��"�̎@A���vy�v��;,
�1.b���;o��CO�>z�w��ZL	��^�g¹U�J�CݵSK���oܧ�\,�`��	:��͡V��I{\�]���'�F�m+�w�WW��v~�'x�G�++�[�p�ᄄ�����X��~;_-�i�dQ�N��D=��b#�S�RW�D>���Iy\>j`pgU�k���:h���]��u��RcU~�}z��>{����[(HJRu���x�ۗY16rh�2�i���^�����4�`�����wp����%��^b�i��r�5�h��^��w�v��6�����b��)����JrVG���0� ������YA��p�2�Jn���p���HW���������#�P�UL�j�f��LR�������w�w����2�'��U<�kr��ģ��U�H�V���o�����H|�>M�֧�f,�mY;����6��{���ы�R��_���+X�3��ZΫ�z�%��o��+�3ڝ��.��Yz<�9����"@������󄈝�ԛ���ڴ`���/�6U�"����ք6�����R$�]T�9�EGMy�q�@������:ǋb�ڞ;>9z��7&;���Z���b�\#��xx��j��SՂ�_����������5Ӱ���qG)�������-m�T(x�q����|X�eo��9���b�߿����5�	�ǽ&��v4ڒ��?�g��
9ޖ�n1X%|%�\��2��1��v��L>.6����B��jށW�D�PK   @jgU�\���	 2	 /   images/ee25a61b-6355-4858-a778-65c1949b8af0.pngt�UX���%XJJzWr����T�fA��A�kY������F$����]��{03�3s0s_��'\UY��޳g��a��Ϟav?{���翝�u_��'u9�g�c4�X%�=��ſ7���Ƶ�i;={F�����o���ٳ�yi�O��δ�M����W{�����^W\Ju����#J�,�u𔔅����%H`r��߫��(2��B9��]��EC2�L���=�N�a�����]���ߜ>>xE�x]٭�=p��	؝�^Z�x^����r3�hIN]���62�/8�]ԥ�>���d75��������fu5������O�����R�{�"l9L��3 �:�q�qU=��MG�/���$��rKKK��G�v��y{�g��Q�{7r9�*v��=޴O�F����[�6�~̎#H$2��AK�ӧ\�E���be5���"������\�A�������r152���u����ճ�\ �v;�'r3�ç�����w諮녫[G�n��
�"O��6.����d��Û2C��&�?.��m�k����?=��ɮ^���o� g4_���	nڿ�S|�-`U��4j���N$g�2����p���� ߱��?bٮMAB$�%w����>/�������}�d���݆�X��Da���f�Ϝ����%M���7vk�}��v��cWB���n΋~w�{PS�/����!�Bx�`��V��ir�|����g֐��ԝ����WFN?*��X�'�-���[��}p\W�˗]��D�27'���ި�?�~�zXZ�����r��6�wH¥!bh��C��)�9v���.;�;�+**�����mB��f��_-c:5�F���� z�}6�j�ZI��~T_R8��R��x"6�&�/��B�g��N�ry��-�O
���^qY�p��c&%\�ҹ붕��ˏڷ�����C��aZ1��̼9�6��CX�><z��<���4�,p���s}�X�y��O+�b�;�dO�m4�khMFf5��>���Vm'V�^>�!d���<O2����z��i�^:F'׫�G�W߀�B�].L��Q�R��UcO}���{g5��5JS��?�c�i����.��͗u���T�kx�{�!,*�"(9���=� �I�u_�i�4�Jlܪ��R�������u�ܘ�H!)E�%l�M=��oz�}��	�,��}�3�Ry�ʫգ]���gL�;�M�ܷ���]�40�����~�F�%?v#?�s�>��Qr��߅�=�<0;�w���e�\I�=@���7�����SΟ&�@�g��єP�����\u�w�"��d�<����讅F��&�,�Wڃ��8xQ՗م��=�Ҙ���0#
�I�4�A(�'��������5Ȱ�����j&��#�%��aN����$��SV�0oor�>���G�.Ϛ�,��a][�X�%Eh��̰�g�<��,6p��EM��.����=�k��!v���O�}��ia��?�sA�j_�"��\�3e=|��X���ə��ijZn{��d�7����A�\fz�i���Ǻ���]OJ?�O0<��T��S�enZ��
	*��~���,I=)�r������L�\��M�+���8��څ� R��֞+ Ϛ��-�����6}��=����W4�Pt�%~`�-��8!�|2}�w߼�3�����:��͌��5v$_i��%6�>glF�BH�Y�1�޺ݳ�PP�څH�=�(X�82����oD�猋m���(�i0-������:?Ξ{R�ܥڡ��|�D���fĊ�6�ڱ=�s��d��2�H�؝0�>o!�a��������s�Y���;��7�p@�.�1����:"�Wu�[1���R9�^���ZEΉ���a���ZDU�z�t�*�}̝�E!�F7���Gqq{�Ț<��䢵��y7Z�V�Z�xA-�U�+��t8	גc�N2����¬QF�\�� ������频�s�l��D�9z@w����ظ)0�[�RFM�aԬ�����37��4��OϟsVL���&7���[w�2�����	�����y��G��Ȍ�d5,lѣ$��=n����n�O��C+�NgK�����|�4�f��=HM���o�[������}6A��?l�Y?���hM�,�iL}��2�G�$$�O���#j��,�����R���j_H�U�FW��-�
Mk���n����{�nw�;>��'�3��ၵj}����Σ~�-������N��^�$z�����$�L�-�m��� =��o������SVVm\`�4C �S�~�I0a��B#jf8���.��u�ޟ/�>�\�^��V�Vq)�ʸ+�sI�m���x[2v��gI�w��k8kH|*�Ќ����p�S8�@�7�&m�;���߆�N~G��o5�7�j?B��6%m~`�ʸ�Dn�<d0�����M��]Σ[�i0G�+m_cp� =7i��� ��������m�x���Z��i�i�%��pX�!xy�L±zg�>Kj����<P�U��Ig���v���´�f��m����z���(���Ρ�o�;R+jb��v�z:�'(�t�I1W����ˈ�A@��0�ژ��5�[d��J$��df O�>u��!r�#����� -���wVp�,�Jڸ%M���e�nr��舆�l�Q��v��h�p��X#�؂�����>U��Ŗﵜ)�n�Y�BF��*�-۫�,�)g��xa�Y˄F�w��f�"i6�ڏ��fp����m"ɢM�E�B����Ȕ6`�p���>~��އ��4�Y-����`��'�*��EK��;�~���CN�c�+f����	��&��u�;5+��?H��cT�h�\�� �11�+�3m-��y@@8mp��%֞�wc���_��IYV:q�������o�UG]��(v���_I�}������Pfl��fv��S��{�d���f�8�Ě����{t�E��A{蓒�'�"�)R\1?��A���ۥq`G��M���,js\���"��W���[Ð�����ň]r����{������Sh��&K�����x�t�%�JL���0ڏ�զ[%��B���[���;2%q��.�*MUwyb�^l�.��g{)q}NM�l��8���*�!�_�O���z���qW\l��(sp~�۽�q=����Ml����o6O_�7��{��#�6���`Ҏ�$��f4@A���ü}KqTQF���3���>�A!y�����5!!��鸉�� ��uv�G#�h���S(�i`��^p�g���#T���YlP%����A4��V{��3VKs���l�i����K43�:�{�z���T��|\�eÛe_=_���x����H{�dg��,�xg��[ؽ;LE��.�����Z��R��c���`�@��:֜�rtE2���h܄g�tޞ���Y��7�V�
qp�M<2�qY8E�0�]̘x٥�G/Ƥ�~�ն���×G�c��uAց�-���]
�ӏ�'�7��F �Dax���g�Ǭ?7��@E�G��Ŗ�R��C�(����MO��=��[m�q���(�6T �|�-_M���"��Vhܠg��
�ᠱ��&ĩ��c0��5n�����箮��_)�OLfP�x9��j����7�Oi�t��u4K����97P�C�Ճϑj9����)�����mY6�����f��g�K����0a���!��%�����fd�ps�̂�MGr:V�M	u����e��֠�˾�Q����ƾ��O��f%Mf���cf����3F�$:Q�X2
z����PA�'������r����Sн�53�_�����Q��;�m�0��(u��3��ܻ�Mo�(��|$�s8�Q�z�h��k�C�(��s��ֿ�U��0VDh�s�F�n0��v�*/+�y=�f8��#�1<n��0a:�	l�bѢ�8YN��8�ފj�<�gܑ�|D5]@P<�����,�Uu�,����R1n�1W}{������C_K<�����E=TK%y��r-Mao�gZ�hSvoʒ�&��HQ�q�t�(L+\�bE�C���{rŁ{�W<*]x��00�����/��)�#7d��&�J����]�਴���|�%��:�ے���Ƀ��T�j�o���#,%&��2�Tu�\b�2��) )I��z0yc�����0���t�m�o��q]�ݭ��T,�z�����P��������
�9r4,y�e���`:f;�
��c`|;X$�b���w�]��ȧmr�S��{�5�v|���YF��Ҭ����Xc	��A����Z�d�qHڰ��O�'�Oɪ'g��������k�Ε 1�G*Î�̨�	�^-@���0��* �9�HG�$�ݼ u-	����/H���(�x�cE���9d�$>3���y[�<��'�![?.�����ڨq�u����v'�-��Z��.���٢�/��{q2�6.l�]>E�˒v]�u�3]�,��#�1F{Y�jY���2=��=���2=K�^��?o�u{�䃕Ь���wd:�������k�z"�z]�wJhۑ��a0�j�t�蛥t�3^�o�LV3��1^%r�֓�-8�A�8W}�TV�M�K}�0x�S��%hQ�`bN����W��Ƞ�7�@�َT������gD���>���":�4̪� �@�S�^��lB���*(ΰGf��fi^���PZ�M�ԗ�!��iDf�a�yRR�gcc5���w��?=��4���}0�q%�
,�JAyB�2���:nu8��4��:؍FZC-�U���~�A�^�O9�\�ܿ���~38'N�MG�q�ۇV�%M�=�2fV�e-/F�s;�t���^h҉Vl��F+v�Y�q:�pJo����Xaps��(��8�z5�D��N!����]���ڛ��~є�W��g���1KӖ���8K��+���f����Ǣ/ͰkV_�s
*?*�%"S��k����`�a���z^���B/�G銥�}�f��[�-4i.lb�&�ֈi�;.z���XkD����o32(#E7�7�r7����w����ĨAnӷݛ�c	>�j��@��AD'W�Xp7���+!�W�G�b��Ӫ(ǈٍ(��f�)L�k�#��&3H!J��/�$M�b�q�LKmА���*��?^�͋������o�;�r��9c]V_S�������0�4��a*�g���V��W�y_��o&�Pd~|Ɗ�����v�8NU�|�ڷ����Hi����&�m�_�$�H^���Q���Y=.�$�b�Ia�L��CBS�K
��,G�p�e;G���x~�On��P��8♂H������}w�STx��s��q��ֱ�VŪ���K�k�֚O+ˬ,G��w�:@�����+h!��"%r2L��T��S��h��4�̲�듥N|m�-dxX"R�-���F�-B搑jiO�RM�j�$.�獵�����t|(R�����`�"]��L�����b��l#= ����C$#4����?���L�#����.'��\��t��#'�E&�$9A:G^��#�Y� �X>V!#;[
&"��ޛ+� ���=e���_�?�'�^C
t �r����J��+<#�>� ��x���Go��oa�s	l��Y��Z�T}�X�?h��`\ؠ����NtL��?�g��L�1YXX[>�Hb�'ȟ�N%h+��s�\�?��ǲ��$��E\�.W�#�Ԇ �NCxqc-p��\J��6A��p�˻z/�{+O�MD�f'53���61�]�'F�.rЫ��4UC%�{����v�V��ZB��G7���,��83�x�e�K̫a�hs�`��t��KvIIs�ofS$q�E�Bf\��S�N���-T���b0Le�'��:6����ɫ��*��</�U<ё|�f�(�詊
�d�ٰĝ��rR�<Y3O�X��^-,��]ܢh�yBB�h���ԏ����g�g�)g�ކ�O���D;����
��O�7Xlb=��n�)��N�J��L4b~/���M�~������ �|���x�W�lQ�7{���+�����$�+��9��(FJ�ʆ��v�X����c�i���:{>I��1�1n�{��K�::�a���7��ԯ��#49�+΃��#_�pu��8d:F�_���z�J�r�&6��^�ACB��JB����TD۝+$J�l����*��c�H�����ʘ�:,i$({��X_� |s(EYt��o	Z�L��^��[^�d�\��>Mp��8�r���8 \b_�X���r�:������L�-�iIEV`*���ϚɳP�����
�x�#8���g�N�/�������L#�P�R��H�ueoe�NZ\�2�de�]6,$�2�FZ��8AݴE'�C��/͎T*-��(�UI�%E����]�u@��;ُ��_��ׂܼl8�uv=�"��<V_���>�j/W��HO�%�ax���Ң+gRK8�8�6I❱L�m��g�@��9�G Y�-oʾ�~#�����c� `/&�W�֫�ȋ̈���MN���q�D$��(k��SL��Ecn e{wzBl��9Wo���ck�jMnH��

��n]~�{�_ؘ.���������=A3A%�{��/��7θ	`��d~�4���Dȭ��U�*�`�pFvdIA����?�`x�텰n�f+�$��
�-~~/ј�1yQB����SJ��S������W��Sc�|���U�;f;~3�擪r~U�����Pc�.'���v�8u�^=B�Fl��4H$ϫ��g��Q>'7�#v��.���Bn�b�爴%�4ы�!	)�oy����½�\!x5�:�
&���)URWA�3o �8�˗���(�Ll:G|�`��gt;ހ����ժ�9e�#rp�X%�w������G,y*�&7Аð˦��i�� �P���˘��m��߫��L����2�������,-a��F)��!i�>0o��,��̀��7.uH�[f��p���0��E2Us
��'�`Ի%?_Te�H4�"�o^]�'��@�b�DJ�^ʍ�;�\�W����9����r)��Z�e��]���)�eeo����0o�7,�)$כ��b>CfЂd��OJ��⃹�Տl�J��ť��P͝
(�J���p�����ܫS��{����ߕPA'6�"ە��7��M¿�NTw����ԯ�4r�z
�r8�W� �Ko
���6ݫ������b^et�</����� ��*�ǌt���\��\s�&�?zA�dB%`5MT�F��Aq���e'��+�)�Dr��䩡�4Rkm����ǏJ�b�!lJ�bÿl>_4�3�X^�s�1�-�ʊ�
��AMQ<k�!} K*P�B�*�SOjTnGt�!��Ϟ��G�Iđ�y�78^ʿ%!ҡ���EϜ�/e��ݜ)�"���MJ&�H3JE'��0/v�Z���T�C�ng�qa��ߓ���4�oޞ��5f�_$�����T�줶�vv�j)��<3٥c/�O�Y[������슯��|&����ٙ�[҇BKg״0�ㄉ^�"6ޙ�ڠU��w7��/��=�3/�_IR���_8�K���_�ä��y�����/L�T��`�t!��QL�0��0�e���h��w;챾�*J�\�jAR��wJ������ng�YT����lgT��:�AĆٶ�*P��=s��?8mD!Hŏ�`�����(�u�d�I
^v��z�t��F]��}���"�ܐ�f�}�Q&���{N�zz�:Д����WdJ�� LDnT+dA���+�6$'��aϗ:�X�\�"7t�FLvۚp-�����'�y�),�l՘QOql/�AM��s0!lm�LVk�zX�Z���aX��:C)n��K�$cK!ԟI�C�}��=�6%ݡ(�֖���3O����9x�!
t}�~d��H��6̈<*���R����
���!I2�Xђ_�J|\�'e�\K��L�qtp{0vĺt��w}4=�(g��iޓ<���l>RQ�Ve�{Dr�Ϗ(1Q2�:��O�e�p����짙���[6,�-)��,�u�G������o�i翳%mǻ"�ĸ��9]����e�G�*�B�Ly.��Χ�Xf�9��XW[n�;pƬ��X.��=��-t5o\ZJ�@|܍�����7�@���2e���-�{�'�U�}��
�n<�i�w$VT����L͋A�0�p��7�PO�XTb�m�5X�A4~3�����+�o���=��`\�P���Zۢ���:��x �uM�[4<�cб�v&\P ����^��Ȣ0��"�)E# E$膿r�<.�+��i8_��Zmƿ���u|�[k�?;����_��9z!�sȠ�����'��t9��xzb\w���%{Ѓ�D��u���˨���@�,��E�T�[��й�wc+}c[��{��4'����?A�%e�>)E�A��up���}_D���#]�n�ѝJDo�?���*�+_��N�jxv���^U��G#ݎLoD]F�6�zl�S���]�q�F���^��L�T�L���!oJx�
J�͘�&I�"�0�]{],��4�cAH�`Z��Y5�C�*_I����J��.wȢ���=��[��-�2���15-7H|���Ԥv�$x���iFhXȉ���)/�9az�
&�}�X˰���"��#��"�H�e��$�в^/ĝ��B/r#ٓ����W
}I��>xy��--��F�<[\�htpvH)��GDz��R^�;,�QV�_�"ܬ$#P�'?���;�tQ%f���#%�lZ@�)���)L�33s>��� I��O��:d����/�TG���W`
�ru��c	|z�y��u˨���K^�\�rt�iE��>������d���̐��.dDN�N&�,���V�nV3��ɫ�R³�b�mT�땤n���ɪ���%p�����.��A�	�""��A#L����/��D�eV���K�Kj�K�2Z��Mdn���l6�tSe�����]zAc���P���S�����{�/��潚�G�\��ý�pχ���b���	{�R����H�U_J:���O��-�~�g���=o#.��p)E��v����Zu�r\�݊
��,���.'���EoA[��z'��ar�u�f�D�~����� _�"+ժ}q�;��ȨX���X*Fߞ��CʃT��zU$�ܻCN� '����9
(��8�����j�b�jJ.ڟlޗ�:d\�v�`>��Ð�~��]�*�����3���\c�>ASZԟ)py`U���g�F:#��F�M��ͥ��`ô���m��NΓZA�,��^�p����� c �nE���²�r�|?��M@j�h�N�\����-3��t�F��Ww�}Iq���#�M����/_���K��0N�o@���f;��1TOa;�H��WP�?�+UY]�3���Riܬ� �tӓn�d撒dx5������UEAb�|�������H\zf�Q�YQ��0����*k�+�9�>��CUV2BA=.95����2$	��w$�+z��W*��`�8r�}Ou�ӒuJre��ɡ>��2�c��{��j�8
U���v����k��B����9��;_�e	>�7~J����%���Q������uf:�y Z����)�}CRG/@k�We:�q􅺿Խ:��m��4ת��?^��O>���+脧K�ۗZ�x�Q*����#�q�2=?�g���J_Bs��Y���_�U�5�%z��9�4K����E%Q�S�_E�_�]�R��4vK���p��	���
������ ��/�f)�/u뢭?+���{̾c�V4֓5��tc0��2&�[םQ��Ow�$��^�" |����8M�P�m�=���-3����M��A*������U����jQo��x����G������g��8$��i+|��Q�.B�����@I�w��!MS����޹��d��Rb$or%�CU>&��z"HF�T�|\T��SO��O'�Z�lN`T,Ga��\(���t����~� ��� ��1*f��jf!�_I��dJ������,qE��O6y5E�/z�H~� ����a����+CB �I Bn���CU<7m�Ǹ)���Y��;{�	�UR1/{bQ,���
�C�,	��uz��\��CF����wӲ�u�(�$9N*��\��Q�eo�X��+''
N�!ה����|�������"�%��0��YLؿ㗖�m�\��C8i�'�U��m�W�2X����ݮs(����\v��N���+������v�o��m	�񏋾(���v]��x�w����  ��V��z����}F�L�~E�G����ҩ������g���1���}y�,����נ���0K���Xb�Ֆ�i�W��W]q�<��^�`+w��'�x�K�+�a�����j�9��2`W���Q.J����p���)@��
ԗ�]6í`l���\t%��o�H���'��B�cƟ�y!�h!ig1|x��o����fm�4��ya�&Yn-���@�JS�������;A�E&��lQ���bb��7I
	UU�`ߣ$~���v���|d��u$��?H�(t˞Gۘ��q�b s���a���.f@3��4�I��-,�k��,��C�%r�3Z5�V �S�^ي�,��X[Ƀ��������>"r{��� )���3���L�*��LR2���<+((`� a>J�'/dYӣ����,�D�S�s�[NOF�����˅~(�/�nB���ޜ�����f�dOj,�#=��(��vH�k%3�fr_��W{�D�A�%§��~��7�k�k�=�or��O�]
�)iҒ�$H*�ߑw�Ăb�gL%�gʆ�� ��*$���h��q����E�_�Va�֑�!�)���?�,F�w��re�x�C�E�sDU�nF�{�գH��{A2G�����=�cc�Þ ���ac�V����Β����̶ Q6��"R���k�����K��}�rʦK��}efÓZ-����"����$W�򚗮�i�:��U�eM��[�$����9V�⟜���љ�e-�%��WG�A E	-�
ZP��5k�	t��v�	U��H���m���r-���_��i��e�����;}�	���|I`�������`>h,�F ��1 �C�'T���,���77�R�O�u?N���JY�.�<3�l&��{w�s�n�,�\�D��O`�wd��,�q��L�(qHl�2�m��Q�6gss�xH|9�]�����r��{"Vn�g�K���y�m���pS3~��(�KoI��l���{�V��»tN St��ֶ�<���M�_p�/O��mk�g�{���4��]������u��ɺB��`"ʨ�1�����C6�ނ`x��FH�j�n��]'/�<8�g�禽���Re]ɛ�e��\ɔ����SD�����q��j����A`R���$���0YU�F��.��з���b��kmKA���Jn�!�o�e �U�x���cO��0<��F��P�ȓꔜ#Y��j�H��혆�,��%Kh>���|ɋV����Bg>$/�vx^mf��O�r��؀&	�؁{��VS�9t���e������Ŵ��r^^����uDz^���h�^�[�Q,����9S��U�����ڛ��'LD�n�JY��1N�5��:����D@��P�ef7�,�R�^�,���,$��G� ��i.ߞ.�;��?5��v�|�+m���5�����!�#۵�sT_l{\�B|��<�~Q�
]�f;����ɾsw�p9�N��r���W'0��j�_4���5dJ��L��k˃Wq�t��(�XS�u?��ѬCzc%=�6����{����x�#���|x 3O�K=�Y^��{xX/��W��sU���dA�l8-�:���mj�����d�+�T�*�H�i��&�ɒ��H�V7��7ՓM%Y;������Z�r=:8gf�<H�Y��� �����VE��hF���������۔9����m�x�x�x���!x��Ne�*y����*P��HC�p�����f J��ƅ{�~�[��>(�����5P�#��0'ף���v��S;�v�9g);���I�㮸z7[�A�<�O�$��].*�Y�x{�hI�e���R�2he㘌B�(
x�zD�]�lM(6�oHҲ�d�����b�zQ�� �z��W��ߏ��M�ch���RQ�^W��g[�����M�[��0e�O��?̮�7闍o����m�˥�ͦiX~3�0h��ZU䜁}Ϗ�`�R�� #�J�,�L�w��]�l�gדNP�k�+z����iϚ_����n���V�r�Ν�$��M�`���c��z7�CN�%hퟅѪ��bh�,��5��o/p`���tA����d�q�~���_�J�%�����}L;_�C��f!��z��)1��{��0؃�����odwA�A%/��3
�H�+��I�~����٭��ǈ�Y�|��u�A����N��4�u�}-��ݭ�Z�3`-���E�7_΁xY����:�Sx�HT�a�����]R�`ycZ4ґ<�F)  Nw{"�dU}�������|{��kǃ+aG/9��B�|��b��%y?����ggGp�r�x�`�F`v�l��*��WɆ���}��1x'�,I�|�����?��Y�z3�d���ٹ D�ݪ��Uw�*W�����K���#��FfC]��J���s֑�un�8Bn�M9�nD�8=�Xc���h���d��% Q���d��_i��I�������k�h�U^��W�O+�u�@ֺX^�*�y��ٿ�{KU<l��	9�IB$�&+�ր�L_�Psȍ��5����	kr���}q%�F���Mh��VGf��v��[�ݲk�.����'�5�8d���"�?/.
h\��1�P��NY�=�e�_U?}=�r�b@~�Η�g��zf��=Z�Sg���z�y������!;�9��u� wVsp;p���.a�@�ɡ����R\�!Жn�G0n��e�)���u�� ��)�B��%�<��`r%;�@��`�h�����XƗt
�1s��0�O�/�(ǨoN�6�v��on%u�DpQ[��4&镶���4R9�戆$�+�$�Gn��d��ř��ɘ����kva��&�HU1�\�gA�b)Y��aZ�����	Y��ӊ)�+�x��s����_	��~�k9s�pu�ue��3��R��� ��B����N�0��M'��£0��_������uB���v}���T���)��A��>��䔨2ô�<���	����ԤY��n�q�/ѐyA����1U���i�*ϭoz"��'��]|��+�8���$�g�q�#K�-�GҜ���~�����XC��&���n�)n�p��85����MԵ�i�Z���*�����0�q:AI_	.I���my�-+mҦ c9�A�f��_��t��vݮh/�3L<~c��g~��Q#�}�@Z+a�ې=_A�Y�jvԶ�p})�r ݄j�P�S�A'�{���
3NЄ�����Bc�9s5��m�m��)I3n:7��=���/AzK䦳��06O &���0Q���/Y�K�)�6օu��L=�e��V>��>���Nh荌J6�y���qq�CsHu;Sm��.���Õ�?�0.��;9ٿy�p'�h+����	�(��v�a+ ���CֲGf~kȮ�;���뢆��pϲ�H
\���D�4�N�ѕMň��um5��k��d�v��j��֊������G\񓅲]�Gf���Qj�DR���(�86B��x�"��QIB���f
�7ڨwx���	��_��5}��d���hp�%,o�S�
�}��{�U��
�a;1����9�~q�uG�u��+޶����oj�ߞ#U�Ij�I�=Q�ï��]{ܒ�-�/��*�)�����X��U	�r7x��1��T^e�4��V:^i���x��c�"����K,�5Xy��sO����%��U�a��<�"��D�S+/��Zy��?�X��:���ʤ�iX�Sއ��+��lE��RnnFJ(�R�KĬ�����[���۷brύ���4:	}�k�YM3~v��";��l�$�k�r�������1ُ�.��m�������6����K��Q�G��b�)\�T8�Y���"�A@~O۱zތ2"��pxݾ����ykD��ɥ�[�O��>���TJ�ا���0מJ��V=��f]d[��깝eJ���;y�9���Y�xz��c�e�aqy1$7a�̣謥�j�{n��C0��؍b~��.Or{^�r���g�	3�!�N:����V�Q��U���p]�tb-�R�V/�vB����`�^�W�&S�D1
Y�F��Y�*��̀C�_�i�g���d�#eܦFm�ѣ?�3�����g�F�j-�s��2��I��$+�L!@�W�KK�6�%&��z�R��0�HH\. �7y{f����Z���l+��)7ԥ�l�Q�Mt��h���m�P#Q� ����'�THE����E� D����E���6֝5v�2w�T?P�Ž��\A���� ��顔a�ܯC�:�`�
sֶ ����h]P��+;�Ԭ�$!*o ��/�^�hA��b�B9����O6ZA��Y�t�g;3�hLTO�䪿��~���>��uj&�УO�P��w1�+�;�1�-[��ۡ�����9B�I�
����9�(X���~T_³.R��]�u%
�T��-�#�iHX�*����W�יz�FTO�l�k7,ϲ�'�Ώ���eNՑ�.&Nz�=x�bl�N@��y�VKl7�%�R��3❪���4�.�j�����yRra��i$zԃT=t��t�F6u�
�nP=՚�<�ӨKkר�~j�Ә�y��*���,t��{�m,m�o^�������sOWo��Y��Y�����O}ywDդ܌f-�������a�6���Xl�Ӏ���Z[P���hsL.MHp=h���O{i����&�;N�iÊ��[�zT��x/FkF�c���O��H-%֘����ؤe�D����爟S���v�93�S�4��/��9|��k�'��c>/]�-�Ŧ�!yo���>�ng���!�_n��D���b�J0������#���'�[4�<Iy�495$7���uC�B���v��fS�?:0���G)�ö����C������%���ߘt�p1IH�xe��ޚ&h��O��)U��#��N'g׷5_�B��t��Q�!6a�$+DEo֗N�W~�R��(�be�|�c�j��߻��+l\&w��XBᜡ*����=�[9�������o�b�w���L��خ�~!2�jF����j��w~]�+D�nX��a"�]��DY���2zD=$��ڮ�6�y��X�,T������;J��#7�|���Y2�T�ZIvN�&��P�����\��H}��R˝C���z��ű��64f��?���/C�;Eᥗ�7|��Ȱ����yڼ�3�G��Z|?k�u��+�l���щ�Ģ-T�d�������[/�����O���RE�]])����T=_t,ؑ�H+�?��F)[A~m�=O�8��j��@��j���35���B�1����M�`1^ w��x�7�4[�5�8�0���+��Q�w�9qOz����p~{sP��Sc@�t�1@*~4Ǘ��;�%�������;	Y3�/va��B:t$��1����1�2;ϛ��_�eo*[��� ��W���&R��3�7�y�=�D����V����b����E>u{wg2����R�:����^7���_�!�5�|��v�3����g팎�rkodݭ�{�sq��fhs�t���KV����#},��<�ti��*$7צ���ZU��B]�"���J���):w5�Y�ܤ{\�I@��&U�6"�\;��$�{����e�ϸ��)�7�$�D�/\S�$�8f��a�o�۝&�r��%r�v�L$�/�8r ��ry��5Aȏ�s�zxvn�D�<I#R��UϦ�b��tHҩ���9@ƿ���iҞ���n�v�u�E$�yƛ�:ڳ����[ܧy$Εi�ʕ����p�EE�w��Q��p�ڴ֫V���5/e)_�Wq�bf����Rp(P-)l
��(��4���)����q�)�-�W�ԃ�zJM��1ӚHo�NK�i %E�[�oD��{[�=�up���%�"�J:)���?��\W
aKʦ�BB�iI�Tȼ�+����3]�iͼ�)�mG�Wq�i-o,ߖai��i��i�i���v�ධ�$R>E��R����{�Rلrل7;�I
���)o,���Ud_$��Z�Zn��H؂ܒqB3Z��H��5'͸]�g��s�K�mc���]����7�ibE)�ӛ��J{m���
\�﹞M�g���F2NhB��6�馂�\O�h��4guۉq�}���.��&�]桱�<�ݾ���f#��z�5�����m�`t��l�cZ�7vo_���gQ�{��7P�q��琗|9	�����_�@^�i2����AA�i���EY�y�f�EI�)�&Fv�A�&GA�9�u	�gqp�ZD�N���Y�@����z<NE߉�:y�O���m�p��y�zzEe��)�ū�$�(	oӕWh_��{�*�*�Z+P�ͨ��^
�������p9EXd���i"�&��}���b�y���ݠX^���9v��ƺ�k����?�ªwR�`Þ�X�{��',��#�mڂ�`ɆmX�yEp�"v�f�޼�6���C̦u�޴36n@ԺM�Z�Qk�!j�6�.݀�%����(,�"l����W#D�'��#x�*�]����.�]��y+1����K���cR�2L��Ʉ���eZ�b��Z���1�Q~��'>�35�/�{r�#b!Yw�F\��%l\B�9t>��й���i�$M8)f�i��9p�נ�p���s)ç�WX�;��j���^�û7D·x]KyUԨP���O᭭�Due)GMU��J�!~#���T�1�߿VB,a-�+ʊ�'o �ΠX���'ذ~��]0`�`t���B�a�1��N��p��?��$��O����<֓��Ҙ�I�(��5&�3n�2��q�>+J�Ȥ5��z�L"a덁�h2�S)�!c`l`��0���1�;�"9��<����ZM��8��؀S>�����`�oF�L�p琢a^S��N~�'=��{� 8R�Mt���1ޖ�oC�g8�1@�) Cd�����sGϑ�<):2t� �	,7�y���Iq���ΔE'��@��A����^��^2��;�)~]=�W�0�B���M9��љ�<��x̎�R5>s�&z��^J]�_*N�PCIaf�����!)�����CA��5���z(��)��(��(Z�(^�)p�Y__�to��͛������eob����K9�Ma�EA�M��� �a E}��L�C��o�\'�������q"oRf�����N}�J��W�~'���ϒwQ2,������<�Of=D�E�u̅��'e�$��Yo;7M6uڹ�m{
m.�7�ew`t�s�/ҟb�i.��P+��R~�R�롄��_�|g��H���
қ)q���Y3�D�0ߊ��J��dX�0�V��ϣ���dX�iE�ii�oMi�z\)|&4��hI�n�v6���i�f�a%���9D\�����千-oTo�����H�걶@s
_3
a��6�D1��(���4��"�=���&LW�T)���DoMqe��Ǡ��2OylBql���=��HSҌ۴�iZ��~�xsԌ���3�9�))����V���{5d!��[zo��T�U��
��M�����ֳ�~�V
oc��Ƌk��=煦�o*��D3�vj��j�u�����K��vc��Ј�md��f\#S�:�ķ�A�v���5
��D��Vf5]�v���H,Z�[7� ��%�PZ��/!?Q$�e�<e�"
IA��/�I^�d?;���'�[����P�.�|/"��d%�� �`}����\<��/�����S��[�C?� t����Q���ӌhl9~?�:��g�Q���W�`�0U�%���Od���(�f�z�u�1ğȰpl��;LB!]�2.�"���T����NV�i2�ST��O����K�{�~<x�w����[�|f,\��Z�Q�W"j�*D���d�jD��%k�t"(���� l�ZS^���XDQ]��K�#x�2�,��2J,�-و�7cڢ��,���9��*�X=\��֞0[W���%}�M�[��s�`�u��p=�w�w�D �9p�jĭ�?������ɬe�),�O�xG/�W�<彈,�{��׈�d	%v�F��
QK	�3�;S��)т�NY�g�.���Jy���˄0L
����ϡ�7.�? o߼���"5x�Zzq���H���4�I9��*CuU���k.�m-EZ$���IOu9�?�CGc����4��n譄x��!��0��c�=0��V�~��OH �
^����^fxb�Cos��0g_w��|�b�����C��Y�R0��8�Y�!��;��K���=)�^TOEkw��>V��=΅8'�^c����my`��r�ڻa��;�s� ���u�N��P粆3!�i��ǹ������?l<&��sl��}B8o������;�%#�ba5u)�Q�(��c1d�\�_4Ő��(z���3у�����o,�c����M䓂��`v����b�8�C(�Fz�*��@������sy�\e�+ס+�S��2���Ѕ�T��,��3)�C)����a��>N���-C}c0z�|��a�a��~0���e����^�0�g������Uc0��{��l��`&�,�m`;MF�i��:⸝��A��.DG
�;��Ni�b��+6�0�TCa�+��aʦ�y-
�I�;p�w��R:uڋ��&���B철!��d9r.�=E�=E\M�8�v�v�:�����9�?����
N���-���/��^�=���֔��{Q��)J���_���S�ZQ��Q=��꽞M�#���!��J�r��k�Y�bU���&�"n�3+ʩ	��0]���\+��8��VQhd%�RLXGP�M��h�%�MH/������-%�;{!�R��u��w���4"�)�:M���6�WA�m̺��@#k.��ޘ���[���0	���u��W��S������k4���hB����Z������i�m��l/.GhlMD�I#N+8����u(��o�8�週�4xz�^����y$6o���GgQQ�9��)�W��x��(��P�~��WP�}�y�P�s�b{��.!�Ź:�)�ɗ	�9�<2�G���H{v��l�3�:J��8��_?�yK"`�e�>6cЛ������s:�{MA�@L[������'���zpP���E9t�b�p���S���Iq}O�.A!�D��la]v-=(��S�_I9ʊ)Ĥ�\R(?��E	�o?x�}'N�瓧���#X��'�޾�6l�l
k��5��՘��Y�KV l���[��e�q��u�Y�1�� ��p�x=�y"E���E���N��L˫��-�H!�������(��)�����9�)��)�k)�k�3k5|f��w�*��F�4�Yk(�k�C���#f%�cV�̈́k�r8�X'ʭ��K>���d�J
�

�2J�28�/�C�2؇.��]F��6�H�X�4A�I/�!�`�6��	���s1~z�8�L����X8M�Iq�
ω�8p���o>~�w��W&������x��դ��g��&�H��<@_񠭭��bA���.ū�
´�
Η+d^���`{x�r�2�8� O�?�ً�i�f,Z�11�8=Ξ�������ic��V62�C��b��#Fٹ`�����c�\V.nĝxOX�zغ�B��7�����o?8������&*<&
�JBl"(T�OC"0%b&�Q��A��E��[����d�_G􂅘�x1f/Y�X��-\��׭���l�F���G��Q�ہ���ٱw?v8�}G�c��c�o� �=�#'N���SjZ8}��\��������8q�>��>�	3�c,��m�-����
Y���Y���>��~ھ>s�G�>��H�a���+�	�O�"�&}7�^~��2��������R L7��!��\=�}��EZ跄y���i�ۇ��^��sэ⨍����`���u�$z.�/�sYJjc��1��'c�G���!v�.l;z?������15v=�Q��L��i�[�<8.�5%v�k��b0`�F��d�9���q�'e���$�?{�< �H�򝁞\^?�9����>]}�����f��H0����z�;������!"���N0ɰ���2�YP�L&�HG
�Nη�W�9$V�a�|}���䳄�Y����m����u�դ\͛�t9�^K4\M������cS/�eD)��C�(	�EI�LK[�OD؄>F�9V2l����/�LW� ��,�r��]���i"���9�؀a�qQb��a�{a|��p�pJ����a��P��cck6ahl+�+��2z�ƶ"�"�ᬓ�	����*�pZ��?>�m��F�*��W���H/o��U����K!�(ä�8
����(�
��Xn�.N`�c��D'�u�@��F��q��r�4�eD ���ڠ�xgt�7�t���8�k)���AE�d<=������p��WP�&|y��,�qV�E�Pv�)���N !���2q�O. /�:J3��U�c5,"��9$=:���"+�
XWI����An�M����-#]������<y3>	='��^�8w6���.���;�Q�����!����#�+�&!������@���5QC��Ŀ*ú�"lI��o�h���kO�ɫ�J�)�E���j���CZz�=�;wcǑcX�c�lي%��`�굘�p1w)"�/DHl�"j�"�T�2�,Z����2{�f-Dd,�(v��,g�5�^��KD��!x�JL��S��ڥx=����� ����9s#<fm��}�z��:�E���5p�Zg!rUN�1b%�u�UÞ�jG��9o'��\	���*��Xkʭu���!���a<�
^�qB�2�Z�1A+4�W�16x�	�5��*h)Y�?}1x���,�2Î��B�	���pL����ϫ��(ïyP(��SzEn����aC֑2�t��-�7<@�TW�M����j�_��o8�P����&	�a:"��)���j=�l!^�L�| !/K������m�v���;�����������a�Vlٺ?n�	�y�m��<;)��4v������={��d/v��{�����p�7l�懓�O����p�\>G�������7.�˸���"��]�?������ً犧$!)i��tE:ҳґ!�P��H�+R�#��-�"��+�FaQ.�H���˵5�܎ܞ܎o��6���M�s��U�}S���
��e�LIƉ3��j�#g�����>M٢��zR0Z[M��#�l�$t��@/OJ��|�6��{!z�|��>��SA!�[Ɠ�R*�e~	ex1z�,Dw�U��Q�9�=摹�8�=����A�f��^/��.by���nҝ��=���|
����K�j<��"J�R
�r�˘w	zQ{؇��how���+6���GH�)DI�;��y�8�!������m퍡��`�8	nAc��V��r��	aX�j�ܺ������[��ry�L�/��'.aҼuh1�]�)���Ɓ��7�\c��u�"L:�S�;Q�;�Ţ#�;Q;S";��^�i^���R$u�\G"�:�ko��B]>�8I<%���ܯ!�xѤ��7�\`Elu��D\C�k���Tl5Lrk������]x���)���uZ�
�m	��sȸږ*#g̣~NW?�7Do�7�r�6h���6~U�����k	�eM 5����f��f������f��f��f�椅UZ�崼�8�Dy�[(�%�mC���\w��?��I�f6�o�r�%��MZ�V�B$Z�-؆��f�-�l���ᦜn�v7K�W�*���X�a%���;���d�,4;ߍ�Q4""�B�13�����BJ/��UD�|Ř�>6ߍ��#���C���A����-����Ǡe�v9b vn���ĳ��s��I�>>���G���,
R��8��n!�b�̸�'����)<�?�{w.���ӻp��.\9�n�ً�KG���Y��U�&�Dv�5�=?��Ǭ?�
2J1I}q��q��n��	�@G[t��C'got���x��ƨIS1c�J;wΟã[7QQ\H	.CY%�2\.�J!�0ɰ��Ê�ꝼuP�u!�$�¿�=��_�5�y�e��Ue%E�(��T�u�{����[زs/6��+؁E��`�����d)B��C0�W�����c��eض}3�e~޻�š�����;���MX�v-/]����E�9�1�c&����yK�׊&ƭ�_�
L���K�"x�L��>���[�^�[�I�go&��:k\(��1��N��뙱�Q����v&�%��Y�i˳.g�)�1뉖fϲ��k��e���.jC�36�a7c3�[6Q�a��l�rMD���%6�k`������D�����;�-U��r��	asp@d����z�)>4B�%��~M�%o-A!n(��+B\S�$�=�L�D|x_����-a�[�N�G0M��@u� c�_3`~�}d�a�5Z�j�yMi�*睢<�WT���BRD�Q^�xR�(&L+d��|��RR&�.�O�g��?[ei�Ygme)^UIX���Q*ˉ��ߔ*޽.�lj����PZ������ć7lME���V��o*��m%>���r��ީ��)��*|��L����vY�����&jJ�$�Ks� �.Vq���H|x�~�� O슦��5���UO���H���x���3C�^h2|
����X
0T�i�Y!�N�����n^�9M1�Z���-p�tc���`��.��ά��E�t\��n�%��1!���Sz<EvM�c]֭Bn�)�t�y��J�;����J��R�r��n�S�u�mă�LT�C<���y�_V��+������s�.b5o�##�1mZ&O
"����܀]�|����+��J��=��TT!��-V8���]��A��;m��F�h��4Vw&��P�5f�����f<�XĖ�+lD�:Q0j^�iH#D���m���+��U2<�j�3�~���o�.�f��q��H����2l�3al���[�\�WW���O�eB
`�kZ�ꥵ,����H�bs:�ɥ%�����Q?�˃[fH�1�oE��(ǲ�ic[�R?�.��O�0�ഌ��2��״Q0[RB[R�Z�����f\(ڎA;�p�Hts�"��b�N�㧣��4�k���&��[M�tڍB�q�D�%a�'\�M�l5&��=c(�l��!����W�;
�걕�[ʽЄ륍�͉�F�C&�L"l�����F��n.C0��7lϷc�8�F�������b�D�y����_��&=���vѯ/,_�����yo����aT��a�Y�<��(͋GZ�%��\F:�8G^��s�W���i��!>�;���6�u�(n�=B�ک�xt��]DFŘr-o��H>���c�>�g�~Ro�HO��cg� `F0�Z�羵�u!�&�3����D�������t�
Nڇ��e�$��2\߱���aKC",ɯ�2R�|�ո��r��^��^�p~v	/����ظe7Vnڎ��R�����1-\�I11�>{f/_�5;®c'q��<z�yOP���iQ��Ź�Q��Y�������q�w?��K�/E��h��`Zh(&Ϛ��9���na�1q�6�.?��G1i��🳃l�_�v�����#<�� �9?Pb��y�V��8Τ0̔��l��n���vm)��"��&b(�,g��6z#lfl`�����Z�[�0�����)lglU�Dm�u����Z�U$��B6c|�&X�p.��]�H�F�*9�r$=t��Vc|�JX-���E��6־a�����i2���BjB{��.�RB���J�n=�о��G�C��Ôa�K)=�%VC�W���6V�$ĂI�?P�?R�߿�PS%����][��o*5�d����UO��2$�l���U��+��PY�2�	�SPV�y�����cHj�\�_�|��)��Hm>��:���,�+jY�|�.Ļ��z*s�tr��\S�8�2�R��u2����L|`(|ʲ �Ө����4�+JcSS��T�g����{y��n��D��C����U�~�S���)�������<���B�!S��Y^;�}��2�DRt{r���]�n�뺐0t[L�]B$$"���Mɲ&�zn7�q7��P=���Δ4�wS��_����s9v粺��\V�mww��t������"!Ӻ����g�������\�uA7kO���"y����e�a*�Be	��k<.�����7�)O�$��\?������3xx�/���(R7QUersU��H�dU��H>��q�&�����==�Nm��6�-�e��	m)���f	�fc�pʰ���5��s5(�(���S(�]A�gy5��F��{q���/[�6�� 2��߰��^���z�<z��M�E.�2�ϛ�,�˰ĩ��tD&�DXɰ��_�e�e��W�Z���h�K)��.ĒO�THX?/�(��Z�V���� -I+�pJh[�nL8:�	E�1��4&�Iۡ�h;�����`��v=���Ж�m>C[�K��eڇq�h3�����" -���	h>p"Z�D�
!�h3Z�a���K�o�G��귌��4��5�W�|s(��Q�"�G��1�*�N$��k.�ߒo�1�\��~���2dZd����X2f:�>䇿�s����M�hڭ?:�쎸Y�xx�8^Qx�<ߋ���Px����Fi�9^*n�$�>r�o!;�E��z5Zr�ed��@j�$<?O!��o�Ń[�6�AB�m<�wOn_E<χn���{����i$>;�$Jw���H}�ى�)���)7�y�f�:X�Gw/����n�i�;�y>�r�6�ڃ{w���p�&��C$4n ���5˴z.�$����5�@�;\'������"l�|u-����.ds�K��:
_�E*%�if!����E~��{�|�6DΝ�Й�)�ማ� ;w����W������(���y�\ʎ\�( ��3N���Ae�|�,Y�/�����d���<	N�^������K�5��-���_�f�Sv�(���S���p�ԺPN�)�NJ~	�4��h���(�n�f�(��R<մ)�����Aa����al��:�����̫؄�a��C���5ƅo���cC�Mg@�Z,7��P�mE�C7`\�Z���c�����a7m>��#�1%���Gq)Ő2��N�5ֆL�K��˸^�7\�eJp?�<�d��,���rk�B]�_�TR0dD��i�p�+Ѯq���+�\A���m9�˹<�-�qRIqf�ե\&�G����Y�{��m~�e�u)�"��G��Ӑ
�1/�����2�����F(�t!o��F��y)˦im^��x�Z����vKۅ�bEu|��G�zz�G����^
��J���ME!^���4�W�~]^��¶���E\��g�\��Y/Dy~*���	�im�����=�M�A������H�������$Óхr�U���Ճ2��k�	m�BW�wv[��zauD�Lb�|"��<4!��ِ�^�d栘���$]�a	��m��&Â�p77
�� B,�R�0q[ƺV�u̳
=ٞ����6 ]����E�*�L%oN���lT�M�������B��<��UXS�����r:�
P�}QV�Û�,�g�0��R,_��$���U�q�E����e|3�҆۶��L��˫��Q~�))	���&���WAv�G	��R0�Q-B�TPr5暐�&ՅS�0ɰ���?&�����[/�2���@�e���H��������e�^s����׺a���	�<�\�:�Ǖ©�I�{`�^�:���G�4M���
�zۀ�~y���g`yMvRg��֟���3<���ȷ\�&�61h���C}����-���v��e�����H4�2ͺY���:ķ�(���M:�c� ��5m��F�Nĵ�N��i���.���m�qB��n�>�=F��'��>#<�o�/z�`�tE���8hz���e(o���:�`Fc;yp�K!nD��^bS��)V�}�MhC"Dx�M�e��I|����f=�P~�&_��0���+��C�-C�t\�6_�sG�>vh�c$Zv鏎�z���w�Aq�-��8��g�P�x
�w!��O(I�����L���Ի��x����=�;�N�уKx��2?��'��q�M�
�3��s��]����p��	ܻq�y���#H|~ ɔ��CH}����#+�:���a�X��s�Z8��5E���ttv	���y�w�.\8��珣��@��ʘ�Ry�+X�A��.�&�Qc���it�Mj�����%X����@~�(�K/G!8���U��zU�4J�KZ���l<uw���?cɖ5�"C	���l�ճ琛������*��B�x�w��*��T�i���PE([��sxI�0|��P�+�2�2��؆(�M��� L��	���p�۩�p_��5�_��Up����R� =�f�Em""�[(�Mʦ��j�F���(�"�&Dt�(��8N�]�1�k1�Ę���2:R�8��X�P�)�Va[Ll5���7�������*~L�&�G�2�X�����Ũ)�0r�XO�+�p�����#7��%��?��ԚD��6^Wu�k��r�3/x'Ea��S��2.X�a�w���<�4!�!2<�Bm�1�2N�5�i�-ɰ�����D�!��%YD��ʲ9�����w,��|xU�G��Gn�z(Ｑ��P[Cj�l���"O5&�����C�t�s;�񟽌ӥ���|s[V�������4! �lѽ� 4j�M�E�V���������+��Ó2<	�g���|�)FIq��Ȭ.�]��V��JϰF��$����2n��aJ~��a�夷�m�B��e��,%���e����d�U�ݤy!���v�p����P�%�(������Ue��<e騨� ���*�'�tn�L�V���,U%��-���b��(E��'��'�����ݔ���B�!���<����G;���mܢ	C�!�!�`y͘��v�v	֑^`ʰ�<��\�.�6H�"��iI�e��RPZ|� i���T�Yc�l�d�+��w��B��(�2�eUϲ�j�"�<Ӳ���Qd-�@n�Ҍ|V�u��2,\_����XC�$�*ZyP��ԃs2^�2�ܪ���^:��U䵡hk=�*��0�O\/���G�sH3�m,��c�K��SZ�W�F��� G���S@$�E,TL	���K��!1�0k��.����|�^��Waն���aݶc�?�{Β����S���®�g���9=G�^ƱWq��U�����q��c\<����츟0�a&z�
F���_��:_�g8._�	�����%ӿ��G�
��p4#cz��"Ī�wt���ǈ�P������(�_Q��$_��(�_����`�hN�f�/��i��=ƢS��ܱF���cQ@.K����Q��0�_D)����P�|I�OSl�!-%	/����[�u�n޸���7M���{�u7T��=��Ei�������v�<��8�������1$<;��g���t/2��Gʣ�N:�k�K9����3n8�ٹ���$4���Vn1rZ���g.c?�E��z4ys�aSr+�I�.µfB�=PW���ߤ�Kq6���P�e��B��qY)�y!�/���"�����8���?��va���q+�-�A�%+��ĉ#�JI@uq���4��#��#���4��o)��osH.���o�)d���𾈢V�i�ć2��'���X�����D��ez8l&��~�L/&����!���NQ��3�Sz�
%Ñ�K/�H�&�uPjE��B�K�l�:�	616�^���1�2+�����J�e�����Qd��u1y��f`���A��<#���ʼ�]MVax Ex�<����c`��t����+��P'����d��j�yUA�����V�d�BVM���S�4�q�"iU�j�~%��k"�yf�[��@�bI<�%1���C���ZI!��M��T��kޜ���z�z_�.Q|xW�d���C�<1�F��D�V}Ъ�h��f��;��/�p'�Y��B;�htu�������ԘWMbE�노�'X�:SZ�.&6��˘�p$�u�q����e��2��P�]�S�W���*t�L�v����a����7����\���FImJIyM���_����,��T�O�Q���|��
R]^̓��x�s�[�1ϫE%(�+@ei9���6����<s?=�����) �<���5]B�V>5,_Y��aʰ�`Wʯ�|
�|�/C�6�w�H;��_`��>tA��63+i�L7�����aK�m��,� �\��5J�?�_�a����/ ���G5�W������eX���\Gӗ��+i�E��"�&!VR\'�Q��J`)�uDq� ������z�!�_��6!i���rZ=�q���������6
-����Ho�L���]��'Ix�"/R3��딐���)�9Ȧ?�� �����M�MAfa��.�,F>�%����*R�((�DnI)��9�_����+TR����YS����)ϝ���W��pZ��E�۫>R�3�z�����w������1a�p4V2�=�&B܈�E��QDdX� �J�����9.�$�a�S�unB	nn���&����s�qh�e(ڵ�A��q~j��Q��e�0e�����1�<���'q��>ܻ)C��ɓ�x��&�޽��Oፏ���{EX!�~���P��2���"ķNP�O"��	��Q��!�>>����</>��G'�xI(�ڏ�1�&<6u��v�S0 p:-���p��n\�|tO�����Rn���K2��jM��?!åu�C!�%�<IE���q3�\����Nb��CX��.�X���s=o.�mZ���/� 7�+��a�-�'��_�Cl���&���o�P�\��]	/0Y�(�DMe.W��[^��GO�a��;0-*~��
�WX4�&��qb\�,�G�*xQ�]#���� �m�:�0�:\B�aA�q�"�&����J�e(�R<.��`+	�%�<}�F��N��j�M���Rd��[Aķ�I�މ�0t�J	\Q��	�6d�'��FY�<ӆ,��	s1�+��ع�8�
�𑲫��!�됞a%�a�a޹��E���ᭌ��@Q�$�����~�k���N�ɰ&¿(�\FC!n�E��W� �/�\���;�˰�+�d�}*)t�OƔI0|�(t�1 m:@�nV���-����NN��.��#e���щ"ܑ'�v�3��0E�m.�C7�ֆ��D�b���X�^����^��&�:�W�0�"ts�;S�)�](��(�=�:������q6�����C�.#��U�(�)#<'VW���h-�Iy`C����g���'�r��?���O���38�
�_�ˋ�S�&e������Q\X�>@T&�d��Eaer��1}l���1 =]�p�q;E����Eb�z��f.��y�8r�i�X�ΎL'F�K]z-A�����/�i��	�IvE���	��~U�M=���2���n~E�)��~	;a����{�e(���A�g���z����+�AZH�0��� �%(M"�ګ���a3���%Ĕ6m�	��8�4��io2���Z��Y�^{6>̄>�Q/�Y�2�@ė\���'���bt z�O��"��R[��/�����|�wL���{Wq����er	�/����q��Y\�s��&�p��A?�GO���{q��^;}���(X{�������ؽo��݉��	�/�w������Lߩ�쾆>�'���hk#�d�6����E��a6ŘP4������6Rp�)f���;J�dިz!6��W:"��_���u�U^�F��	��c��x��&���Eo���H4����v~}�ӏk��t����p
��E�(}~�b|y�O���}�x�G\�x��z���^�&��)�J�Mܥ߹wM!���wX���y��G)���{���������3x�����F�Sxyw/�BQ�U�g]Gv�:���\�.�hb獦Γ��c
���3zv�	�N�Á���2)A	m-V�\�m5�y^�'�p	�+^,XN�R�����/`큟���A,ٹ�+Vb��و�={���G�P^���<\�M΁���{y���_R

��o(�J	����@ixG�zS|W���"��E���72�� Y�S�Ƀ�c�?��^�ap�	�h8.�۴�pZ	�Е�]���`����*�d�o�
�:%���Wdv�������RxEz�ȯ���`����1j�*�]m�q�D��z�s~��3J�p�Z
�9C'hB�3d�����c(EXN���p��|�,
�K(d5x])o/��oQ�x+�)Ub���{�+��]5���R��y�p)މ�P��S�D�]�el��P�TS=�&T�p=��e��H��7"��;ʰ.�ꄸ�2L�[<4�!Fٶ��?�(2\����2|��`����o�u�6]ƢuW;4��l�a���pg�3<�yq�������5��z�M��	qg�Ko��1��
"�j��mLC~�W7$Bz��I!&.�+8s�D�X���\�a�K1�'���1�k:�l�)�9�zW����ʳ��Q��J*j����K�oa3o��-6ѳbZp4\�am�	�	�����(�C�¾�gp��C$�����2���yú�X_^1�إ+�=�ƻb��t���>^���Ͷ�V7J蝖����H�w\�Δ�N"�&dZĸ=�X�0{h8BdT�WG>�;߄��]M6��ח93NG� �hr��(քW�B�Q��e�.�!��A��e���@�������d��#lQ�Ik�m�>��ɰ.��>�P�\`m���iy��z�L�l����(D3�8
J�ghc "�F��4h㊛�+y0��5���&��U�ѵ
���~B#�J���H�S�wD^��X�2�o�I���Z�xK�(��K��L�X��퇁����9dW�ֽ;��1.�VpvG���nOO[8;��<��y4;���'NN#��2�NC?���r�e���0w���������0
w7+�8��Ё}ѭS�۹���Kȧ�l�w�����0o���v!�5��6�mI�'M)��	�1MhJ�m�}֘��Q��2,���Kl�a5,B�ɰ�;L�������Q�YgZ���F=�8�/;�D��}ѴySx�����c�M���gQ�t�Ov���!�˹����{n+��ڊ�'~ĥs�p��)ܺ}��\����p��U*D�%��U�L���2d�&���O!~�G��߿s�1y��"�_��;����A��q�]i�gP�Oюߋи�h5z$�������=���#'N=۰��!��y�=��Wt�[��F-���ϑ�bEQq!�XiQU5�<�C/b%x���`�F,޶Sbf`Jx�mZ��/�F�v�K�j�H:�8(���M���"����Q[����t���C�*��n��!y}�>��qE�����M?n����8;abT,l����?Γ�a�b�N�w�������K	y��5��*	^K���N]e&����� ׋��)+1r�J-�T)�	����:#��6��d׀���@�b�,F�k2|��K�_��-��w-���{렔����b�T>~�U��2�k�^ז�FdZ	�eD��dX�pC��k�[*48�$�g��C�WS�5��y QN��,�>g����kk4~-o�0���c0!�G�p���Ц�@��8�;Z���j����?t����&���lt$�)J�]硧�� �]�P6�RvE�)���� R@��1�W>!�տ�V'�L�u~���K�m�٦Δ��Nl�s�/�9���R�Y�q�����t�����p��ST�ơ�]1J�QY���]��g�`F�B8��b�+�4���b�'j�^�b�(G���°�n9��ǹa��/\}��hՏ�x�	���Q�?�����(Byu9��
���i�MC/���K x��g�z�D/�OO�p����V*!��]����~'�2�z��4�<���jPh�^%����V�d�M��К����nf�r�ɰeZ��f�ѿ��e�OeX����i.�iAt��aK�A�էU��M��E�gӃ~�_�/=��2L(�z�pKN��b��,ǰ5�����f;H+Ƴ��e�InA�jN�m:&��F����4֡�	M�BT�p�	�̚�M�up���2��6��A�#L�3�ha�h��F��r�?ڎ��n��1�! ?�;�R��?~{wD�_��~4��'aŢ�غ~1�mX����b��9ظ&���a�9ز>?l��7�Ǿ�˱o�rػ�����+p��J=�'�n������?�ʅ�w����vq/Nنi�<ѪYc��݇vU���erD�1��n�.<�:�����f&�!�)��Hno����>���Ɣ��F��ۑ�2��K��WuBl�V�GP�5�dxd�iZ�����8�O���.#Ѫko�j�s� 7�r�� ���5�g�?ێי��&���nĩ=Kp��z�?�W.T2|��yܼu�R|�\��_����{wn�۔�����=��{�(·�5<���������s�N!����i�Q�_$�s��z��8���7:xN���'�x��~v?�{v�}��2,o���]VU֠JdX�X��)�e��bRD
�W��*����!�X���^lؿ�2�ѫ�`��%�	����q��T�g*��8�$Q�֦�� �RO�*EMI>
�S����l����Ӹ{��>�������JFiq/�"�r�yi��d�=��Uj���j$�>g;���	n�S`���J����2<>x)ƅ.��`D)��N�EW�a�	9EX�$ׄ.�a��q���iʰ��`�'#7��j��_CdW�@���C��	a���7�]���?{��EQI�z ������j2,c� �x� O�EIqE�������"������o�a�����?A�U��I�߿Ӷ������Q^MW]Q�d���Ç�@��ТM4m;�ێ�wm������:9��)�_�@њ����6v1[�a��s,e8�2,o�0�X�a�S���+D���`�t�{-��ϐ8��5��Gx�cr�����RTr۔���7}�e�x���v�;��<x�����ago�O	ǌ9��h%f-\�y+�c��M�^��]1�u+�Ia돡V>���_Anq-%�7��E~aʪ+Q\S�����uJ���C?
qo�i������vK��nY�����a��d����&�J&u>�6҂�[H/�g�,��h��F�pk�Q�)­m)���V�ƖƖvJ[�� ф�*XS*��iA)��ZQ�[�6�a�����$XBK+.�bܚum؆6lK[�4��=廃od�WǙ<>x�;Fs�G��H�Q�	�>8�>:��h4/��!I��ԛ$(z��*�y��t�LLe:�F1Y�z�N���x|�r�R�G���Dt�c��e������ӧѯ['���?lX����P�����,�%�8�Jr�,�	��y3[�����	�.y�W�/Q[ƐԔ>CY����(|ȴ�x]�׾D��|�����9�7�l���hѲVo؈���X�e7��o��D�����_���>�����鋿���_{�⫾���~8���#Y�o*F����0|7<�FF�;��(2ze���<EX0ȰE��A���GO���񗮶�c�Q�����U[t��ǏmCM�Sd%G^�>�>ߊ��ہ���|�w�ŉ����͸|v7n\=FW;�7�S8/R�/k��X�i��br�6������{��q��
�S��#N�C��xz�ޢ_G���H�?���� #�2�(�i�p�Ə�a�f�G�F���'���k�7�����G�k�.\�z��{��d����э��{�E�KPJ	.-/ ����������a��>�߻K�m��U�1=&��.Ƶ�PY��=E�6��He8�׃$ƥ���լ� ��	H|��r�q��\;��w�_<Fr���{F!~����fgP��Im��1/��{\����T�P�k8��y<��]#����u�=�a����1�Z��e����5}�I�-ȰIfE�GLYa]��!ov���KD�r��ȰӍC'�^ʰ�,�p��>p�3\R��;������o_���2,����w���}4}"�M��K�y7VB�2�STe_$X��`�a%�&�[)>+�
��Y��E���(�J�"������FF{xN~M��,��c�������KW�p�h�j O���u���v���;��S��4��ټ���l/_F���nq��<�B<���dXdV��:�&��sc�E��3���"�!|`��鈡@������tz�����e�t�9��_���|YM	
�3�����nb��Ű�s���v�w�����-^����[��49IY�H��Gfq)R�����}��`�ƟY�b�{�b�8/�醱��1o�F�g$��j����KT�}��w�p��-��E���z�zS�'�������k��~%�9,�,�s;�BLևI��7J4� �#����a���e2��{eء!��S�f�!��<��ـȰ���I�E@5�h�D2.����|���N%��xt�
V4b���(6�u4F8=*M��L�|�Xv�t42U��`"�	=�.}�|7T��F�&�a���Pa"�����ˁ~�/��ᇿ$�%o����7�)y�zp�Vn����/��\
.�Y�� '�H��b��2Ȇ��.h���}��u�^��k0�mفܼ"\<w�ƈ�p���eg�UQ*)��/�$�"�}�ě���(ϡ���˲g�Aa�MJ�r��P]�|9wP�q9I���4�2�"3��B��ߢS��ز�G<IIǬ�Шk�G�^�K�q�SG'��;�\i�ok���֖��?:9�/=���	h12m��ƃ70�Fp�C�a�h<"
��w#g4�aR��A�ᯅ12Ԃ�Шi�n���a��n$��<߶j	{��HN����H{~%�G��p#ʒv�c�E$^ێ#[g���ո|�G\=�7������(�ʰ����'��߿M�%2|O��E�{Hz����Ž�xps��NN<���x��'��q��h9�m]���-��}�<3�O���q��Y5L�>�d�� Ö{��[�a�N�����߲
ʯN9巔P�(�%�y$��N�7�q��3��a'oކ����bfΟ���`?��E�)2ٔ�t��M�%�N����S�7���۪\$<���'�����~�ܾ�܀�����T�g�� y�g��HEjJ"�R�������BJ��e}�?�@u>�ʲ(E�L�yS�GO�"4"�F����D�L�8�`��0�a+0>�"�B��(ʰ�eXʠ��2�A�5	���	%ú,ו3�$x�u%��$����߅A�9-qj\�_Lq�_��޳0�2���/�q��uL�2!S�x��&�޿��j
��J�9%5Ueعc+ڷo��a��y��XҪ���R���@y��Cy��5��(ÿ�>�彈��������L*�+!�ca%Âb��
��G��B�`B}nY�������
k2Ly~U��T��M�k�
q��A���c�С��k �t�o��ş��-F�����������2x"k6eD~⍦S�]cч��ez�Ģ��6A��G� ��|5�w�ɳ��t�5֖��c!,C�`t�N��i��9MA��M�y�9<O�A����exϓkvi���~��1�ʑ8`¤ ��c7={IQ�C~��"�F��w���J%o�*��K��x��ǓrZQ$f����5�}0`�=\='cÆ����r���0�� �?�WB~3���=���w r�2�L����sЃ��j�t���vuX�=4G9�$o���wSX�3Nd����u��7D�D��Q25Z�\+֣q��OEXZC���~mL����t�ՇX�(���-laӼ�_]�"�@�%�ݺiӼ�O/o7���p��\�ɠ���w�R��P�E`�8��7��8���E�ӏ��߃i��j�/�c:�i_�'L_�������<��|?�io^�koʨ�/9/|%ӽ��^��K/7�Q��?0�CON+��X���3��5@�\��]������GgG.���v��]��u�q���X���h|�s<t�7}m���n��>�(�6���Əg��G��h��
�G:��P4�3
M�A��c��9�;�F�����O{QQ]���b��Qگ?�9���T
�C��CA2�6�JL���DY�-%_CA�U�2�)����K����9}��wQ�uyI��?;�,�pE�-f\Ū%�hE�ܥ=��ځǩ�[�	m�l��t��W](�
n���kg{b��t��v�����>�@oW|?d"Z�
E�ah64͆E���(M���X^��?DG�_�F����`��I�|7�7R#���^���c�����m�!hԺV��EA�=�f\@~�I�R���Fe�)|Ƚ��;cqr�\�_ޅ����+�p������%ܸ���$��2|��$wq�V�Bz��)����=$>����xd�������ѭHO<��HI>���K����݋7cy�����'l�±��1�=�3.\>���5x��-*y����%���Wa��a�e�� �u��a��G7HY%%��L*D�K�8:y�P��py6J���'���`�fĮZ��+V#:n"���i���I6*�2�NJ�%Q��K��~�7U/ԧ���]�_��Ӈp��<�w��I(�IGYA6�U�ϕ�B�pA^�ss������4���q:e�ŪWQ����2̶�{]���l|x'Ot�c��	[W{�p l�b�o8�B��&�DiV�}�EX߫ɰ.�����X�<Y$X��'�2-q�A������ga�G4F���/G�\����лw7�;N��q��E|�vJ���Q(/-Ħ�kи�W���?`��
�6tB�����(&J�E~��3D����e���_\�͇E���p=��0o���뷑��S�u���}����ĉ��.������j�>}��C��hٮ�����7��*��R����d���(���(ó�[d�r,2�Mz|M�5��Y�������6��Q�͐e��R�9�I��AG�@��^������Gq�rZ�Y��b�8�����(�y.��%��}� \|)�CG���q��⥫��+�ɶ��ߠ�U-*j*QRY��"�E(�.Aim)J��������b��\�VP�{�^`��S��E�A���=3c���RN�<��D,�(�P��ldf%��'�r�1v����5�>.}e�3ŵ3e����2<�ӟ�pC�,���ұ$�y�0�a"��9L�YB����,˰&���0ʰ.�����a���f��f:��B%�z^)'��7�mBZ�r=l�5�A{�l�A��=��߻��O�(��(���SOG�����ۑ�ꊯ(�_p���I_N�u����>��j|E�d�,�ÿ2�_(U����H����*�F������2��>.��e����\��Y�_��/�P��,뉯{��P�u��Ky'���(�͆�;����C�?���7m��#Ŷ�h7t�F�F��j���?7ŗ��ۮ��-��	������-���n�j���V�o���uS|դ�l��ZuDӶ�0p�h��{ ���p�*���}�����(���T�n�e
�yJ�e�Rl����ȸ����(L���k(I�,�b�p~�e�8�髨Σgޤ _�8_@ֳS�(Ϲ���kX�0�}�G���{@��WSҿ���y�.c������_;R~;��V�Bn���h
�X�^b�C[��M��0����&�F#�2nXz|��ay��H��&�"��t�ƣC�aO����a4��8�;����+P\t9�gyq�O#��QT�2��l���=���n�?�����K�p��Yܸq��CIq�7���6EX��.e�.��#���}%�����L����1� 2��#�B��}��|��F�~}x�0��%ʰ�;�B>��G���s��k�W�S�+�^+Vo��e���dX	���-�(*�!Y$�qj �E�t��U�X���
GFb֬H\��y�3y�:����7��y�)C	�*}�|ޙ��:���7��q��^n�(�Ϥ(��PQ���"��8/�����"ٔa���!����L�DNV�7��@��f-�RPBI�����%x��BB'c��Ѱ������	�u�"%ã�SR)���'� �u2��6�K�q�DñÖdx���&8m�aW	-I�o���^ay[�
X���s0�{�;O�8��8x�"�n�H�k�=|0Ο>��C��7:DX�TP̛��k���o��?����e��o�����_cY#��'�e��+ٯ�����?K���aM����N��%�˻�q��~�8��f��w�m{�eǡh�y���d�#e�ex�$
����.
�(��#��y&��ȃ^����_�῝_�a%�2��Q�7��C$�O���[<��D�_T�����;���*JyL�T��'����;��S�s�`�:�a�5���^��W�D�V����߾f('�J�`+PYS���pM1
�
QT]�R��
�+�F9��^4&OB�c`e�M�w#=#o޽�	]~�+Ļw<g���I�����6�@o�0tN����o/�R���Y�mez+����Z�����&��#��as�9�����dx^����v�9-ol�7�&�/|�?�����ǿP��H��9u�7�\�m74@i��F�)��F����%ߐ���SV�)�����=E�bm@�$_�e^���p������Qe�����yc��x��{��{��A���qwwwK�wwh�qh��$�<������}窪P�ݽ��}�}w3�w��U�R�V������D?yT�C�C
ͿA�P�[�6!l%�F��G�����."�-�?4�`��|�c��z�f��ƎPh =;/>f��G�V���`b���O8�GoM��� �9�c&CU���׆_�X��c/��;���������0��;��1q�������.^8���b��n$n
n�&�:���o���׈n�7?�p�B8�\��u��\M�mb�6�l_}]m�����~�;Y�ִpDO;~_D>�W�/��$*&����NLdS�2�!�}�b�`���,��ڎӉ��p��YPíy�f��f��"���-�_�p?�����灾�l�kf�Sg����1�r/�1|��.�9����pz�,\=�S!��.$_<����p��e��aq_��l��-��{� &����`DW	�:L3�G��{i�.μ�W���ɽ���5�f&!O,s�`�ֵ0r$�<0$`��f��Y��{���9���/���h�����b|���;1\���A6-��w0u�jLZ�ӗ�BܬY���f��C77��#|_�㍘MN`8�-(�IE��K�vy/�]��6�ѝ$Te�����$��PM W����Dp)�������DqNv.2^g";3S�:!`�����ɨ����|k��_it�q3�:f:�&/��tѲK�J�#F���0�)����eV��by�-��Áq8q%��'#8z��y����1���|<p+%Yj��UL�\^Z��Z�^��G�nƲ��V���Z45T{J��C�#��0L�1i="N���Q��0�{0�ʇx?9�Ť
�#�D�p��3�n03��P�Ԇ�A�2��� ���a���H����0bb�0�ѻXB�U�<.�Ü�M�8|y'���m��=G.^�>=rZ;���4�C]U-˗&��v�'�(/gE���^�����a��G_?,Y��2r��w{�;TUգ���oM=O4��u�emC-�Y�T6����eU}!JYV6vT�-�Q�Z����E[{���W��AaQ	�v��}X��EC}1�]���*TտEa5���]x�Y��0 ��C��A���p'�%�A~��ßF��|NG�0+0���"ð��@a��!Ë�a�J��|,���m��o ����g#1�p$��)p]cГ��eADZ�E�1�(�7��Al��!�p T-�J̪T"�Į�V�*jL�׏�c@��7��Z���۽�>�\��kC��6!R�XC��^va�iο�]6�')�{E�p/�H	j"�kEoS��L���l��6��ן40*n)��=��9��]U:F��s_-���a�����Q�
�����Y�X�c?FM���'�]Ռc�c���x]P���߂��\I������%���X���r\�q�^�%�R�X����;��������n��P`8E�p�ɿ)E �<S�7U�Gc�=�����_E�d�;EM�=�\9���pp�ñs�Q�����'%��t���H��M�q��Xf4F�R��~�?�1���;#~g�#��h;�|S��2C�/��.�'���׋(�V�Þs:1��<���H|?�*z�`+��X !q���ى�L�QB�=IDSF*��@➅�vb]?��IGp;���N�]�gzo޺���q���߼%G1#f��'a��ⴻ��X��1|�轋gi��!�p1���9<INAn�U��y�w���-0ww�@gO���apH�A�1{.�Ƒ���r	M�Mb�_�*����MB	�]�E��n5�pU]9*k��|T���rʼ�Ro#n�*L^��f��셋X�H�I��'�|B)����w�x�N�f���!n];�K��ġq��OH�r��h�ACe)�)�RUZ�J���-/���rY\T���"������!''���Q\�C|D���^�P�V# ��^~�<��"hb<ܣg�+��N��֟��9�l,`�x������!������ף�E�k�"���H�~G���?Ùq��E0D��XB�q"�]F-�	u1l}��?2w�����302փ�����X\Ն��
VH�	.ּj���x|�Ua��E���?�g�o�t�\	��"�&Ѫ����*Ɉe�'���p~+"��Ǥu$����Rd�?Ê~���.y߹d�]d("��X�0\��\J�tcG������VF3t�`c_��v�7��!a�A?�'�X����bX���u�f6,%/�Y�b���+����1��+�L��(@���ax%z�C/p
~<Ó&���xL�Ԣ�����A]e*	�ں&�U�}�������e��4�����PZ%7Է1��j-+��!&m����O�b �7@s�;���w-�}��!���vC;+�m�m����W����3&Ϟ�DG�b��<>��P[Sʂ��P�@U+�p�S�C�s��a=Bnx��R	���=�@+Og�R�����,��|-��(+B�����V�A���Y*!X�В�D��0,��B ؏�[ 1��W<z�₱����J����a4zیFwⲧ�@�H���hy�oEG@�(U��q�i;ZvU$8FI�r��&����8F�����'��#��J`�ܼ���>#��)j.Q򌂚����g���A�hf,�:�C?����s��a<�s��J5F�.j����e ��=��AŃ<!�&,�]a������j
ڑSӌI7p��KdV4 �9|1��]��;Op�UJ� ���.^���)x���
��&^A��ش�b�GO����7�Ν���h��Ae�=b8Y�?�pC�m	�"�|�:G$�y7$�]ů���Xn(}�oK��$�LBy�ԕ�G~�]�\>�t���G��E�C��C�8'V�1C�fb����
�4�������a��,߱���e�H6c��f4c��xh�O�.���>}<���5]���p�}��d�:,�O�}�E���Ps�,u��n�zgt,��X���������$���E�Ӌ�����ckp��F<La��)ܹq�n\��Iܸ�$�oRo$���+�I��n� �o
,�\޾�B_'�Sq��Mܻ#��C�1Q�4�se�QH ��Z��#O���4�I8��@t�g0���@�@xL��݉�:[��ۚ%74��A�a�������W9
�Ê���;1\$�p��m�w��Ո��c���ڟ7��,�3�塝�mkΔ0����=�k~)��,���K�o�r�=��Oo�h��DmY1���J�T�.%�('|�KJ�a������_�������͖0���
�����y	��w4����V/�1l��q3��
�S��y�z���!���8e���cXq_b�D,os�)���5+��~7}G��|N�XB�O2 3������>İ��F����W�w�(�����|<\�x�+-�S�O�xӆ��j��V�`������D���e-�-_n�aV�@9X�	QD��@n�]�x^��31,��.y�e��*����3�&F��}1���(�6U �5���do3	������.���x��<����l9	&�K�{-�5����#��a�"؍\
�ȥ0!0,kV�
�]1l,�v��Ċti)��+0�c2�f�G��i��*�bj��
4VW�n"n�V.o�=Ąi�1��11�r�'Վw,lߢ��VZOt�ho��}ʟD;��&�|���#�\��kW��֝�x�Y�V�C�qQ]-j���p[�M54~��M�`c�++';~�8+7|U��_��r�[�P\݄��\Q����@�{�?
�"3��j�h��/���R�J�#d^&_�0,AX��")�b�:�1�w�Ά6���<=����:Xj��n������6�>q�fEL�}:�E�f0�{<�O�@��\2nb��*����!ޓ1�7N�`�8���M�hxN$�p?p�� ��P��F]���:��+2�єBt��!�D�����j������4W�0fx�\�Ά~�L����2C�Ca��[��y���Ιf�5'�\G~]3-�c��^c���9�T7�1�?:���"9����J�:r�#� $j�=���Zܺ�Sg���m�Q���W��u�ײ�G;d��0��p�Te_C��k�M���2�kr	a�N_'����˨���o��@t��aX����2⬡�`˾��K����E��.����]W_�E�(���\ay�a%i��Um�>zπ&A���V���"���gs��ܛǊ?TeU��Pw�w�:��N1G���D1�����	�Uąvn���e:+K��b6�vE�a������wΰ����s�}z�>��g�И~��IW�����~~�_:��+'q5��^M��kq�༞J 3)����T�85�(&��u��ܒa���� ���GwoĢ��&J��Sd-��N�0�N�&a8?/GN�����CX6��q�)����I�8ǿ�@o{+�~C�EB���v���3+"AX1�Z���#�y�Q`��=LY�F����3�aߑ�hj�!�
%������|(Fi�]$�݂�[�cזؽm)R�����pn��X�B�R
!,��E�.--V�p1\�"q!]a>1�����x��	
�3x+�	L�Wㄝ�'E���x%��8��-z*<&-��BX�BYy�8�UB�(!�,�����=0̌�z��Xn�v���a�	�1e=|F����E���
�w�� M�������wnC�cQ^6J
r�����O�2R�A>6f������za�Eā'�1��?��;����{�p9��� ��akb���P� g���Ew�P>
,&��}!\�A�i�<ĳa26��`:��%0I�F�|	�"/� Vj%�@���0~�~<�dYF����4����lkl@sc+޼��Ҋ�ް6n�p��Ů��PT[���VT�֡����ϋrR��I ^�f;F��h�"���?8�13p21	�5u�a�X�Lp���kiC=놦�a�����9 6v�����\b�=�����5��7�5��gi��foL�Y�b��������Ŀ0� 1�|�c7	�-���������03H�'�3��!�]&�b��B8�l��s����0'"C�K}��.�><p�Խhh��k��
�ep��I�cP�)�\O�&CT�u��K��mM>&H�*��5b=m�N����.8b�_i�~�`2��� �2r|�c�]FNY��f���%�5�2}&��&�G#��s�7a�¥�;D�vΘ�f��=ż�ah��I3p�i
�[�n�1��0c+L��I�\�/�#j�Dlپ��h�ل$��Ga˖ͨ�(@]e�E7	e�Va�����8� NE]��"As}ಌ$��_&~S$�����RQN������I4��-��M���=��مgyX�� �=�`�?
�Ӥ
��Md�lt�q�Ŵ�3���^.��M���?Yx�?-=�g3Ot7!�Ņ���Pu�5�IPu��~�q�!�E����b�51611��8}�#�m�;�sA�oâe8/�,r�E��S�&��SQ�=�W�mB��HI<�k�O��q59�W���̥O ,��qRgR�'�f�U�u�6A|��M�%��	߻��D�k�q�M����b�q�)d��)\� /�v��7h8x�����kl��>����5��A�.��F�gX�2�(��?�L]]j��:���+a��Pj�I�I/^��	񈙻�ΞBYY��ޒE����1���~���?�ı��q|�Z�>��^���Z�Ũ lkkP!,O�!\���"�*L�"����!�3��Wx��1^�x���,�\`�ZB�7��C�vdf�cLl,܂#�=6�#��9e%go��t�_�4���WX�_Y�c��#n+��6
`�(0L�vv������f8� ��q���h�=zC�G�o[��y�v��ɸ���6lE55��{����V.Gr�E$_IDJ�%�;uG��m���.%`��p��VWU���K��]�4%�h!�#1�������b�k��}'���ѹ_~+�+�t�,ƍI;������_�ZÝ���>�}�K'}��C�b<��A�!�m'��u*]�C�ut]���>z>�0���|�r��R:,�O�Vc���R��/�b�#������RL�x�b��]�SR#a8���'����ڸ_ޣ��{�����7�����ˑږ&�3bԚRԋa���v��a���byaa�%u+1�t��k ��`f�� ��F`Î�x�_�Z·��=�Ob��x�W6���s02���(��>K|נ�UL`S�򷌀�C��
�����R�'� �?���~-_F�o�ß��c��`E��a%ߘ�]�}~;G��
k�����ۚ�6!�A�j	 ��Űi����#r�� �<=,G�;�@%��0�����,`�	_���2	`�~�$(!�08t��}��f�.��-����30ZA�).�c�b}�Z����c"����5�ǉ5y֊X+?��߭�o��b�Cg}�а	��s0��8�&�bj��7�|5�&fp����T�*)���`��}c6�ala��+���b��x�]��Wo��'�a�PC[����6Nغs��[��_D���M?�� 5�QUt�����EB\<�h�-��)�n�a�ʜ����E2W�Ƞ��,����ji�m̛;�r����2K7�/��a��diim?V*|gK��h�2~3��7�>qq4�b����^���~0�\S�%uUQs�U1f�r밧�*İ
1ܛ��Ep�&�{�i�Y��1�-"�c��x�}�0|��iV��!7�4r^A���~����kL
%����zn�R��N�E�"2o�&��5a�EDK��k�ۗ;s-�0NI�k���p�F
n޼Τ▄�҄bJ�\>����������i"��u*
2��~���7AϑǏ�+#a2f*p��m'���tbh51�����������J�^���%w^�� \�B���d*:#f�k�	�21<z�|����e�6���4���G�xC�k�!��%�ԿBR�N�۱I�wb��Ÿ�<�	���b�T�����Ly9����2	�e��eI��#\�����19�+�F^^r�2��� ~!͒V���Z݉/Y�b�4�DqI!�o�sG78���G��w�����7Ó'�7��-���."Jv�Y�ޟ��3�1a,�X	ò�~d�"Xb�+���l��8a+�6�7�f�=��y�i��Eo��u��ac� ��# d&�§�r�#�Z�*}4����� L�4�Y�K�p���Yb�ԉ#8w�8Ο9�@?o��?�'��˿c����^[�_[X��c0�5�u��������GcXl���Mn��%��EL7�V�4P��P�4F�������[�� t(K���`�~�ܡa�av!P�u���)���'���z�h�]�ȕ��[�6#lú �k�"�������7�s�o�Y��h�Ђʺ���&��C44���3p��G�Ѭ��@e[*Y����KO4TW���	/��v��L���_FDMƢkp�������NL�O���;d,��G��6�����e(,kByU3�J�Y���b�����-Ĝ�a`�鳗����nBs����R����{��nE̪]0��%r�K �aX,�{0�����+���=��9E���z?��B��~�2˦f�E6��b��`&�����k�����"���A(kp{�ģ�:�_����@"d��l�5����(6�u���M(��ݠXD̀1�T��i��L�����1�F�X[�K�?�����$p���u����<��$�΃��l���"���6��tF�/�ӈ�g}9~3�)��h�dT}�A�{�4-����������0�(�,�ƭ������JX�;a�p}�F��s"�i^�?z���w�90��jSٻ�����p��;ϲ���շ�ޓ�\�߮�҃���l߇��z����o ��MFV�S�6�4�6ʉ�J%����7�Vaq]=!�h��-͸����NFM�u	����\��"1|��ɨ+��{�ObD�t��hېYR����H�n�9��e0�3��7����lzڍ!N'B�+�">���4~obj�I��8��C��8=LB��:J�N�j�4�tO����NP�D?bXb�i��t"xzz�BV�z{)a�i2Ԭ��{��uA�Al0���Ȧ��!��a~�C��8���D�r��<�3Nm_���"��$'�@��3�|��\I���$_��L�E.�/I��d�R�+L2��\C����:RS�Xt��v�"RSp�v"se��2O�Fn�5Ԕ>A��|z�b�/;�ejmWV0Cy칅aX`<'�c��#8y��\���ƺ��I�����߮Q�p,���&���@WCW�
�H�$�R�y���1|�V�̘����v�6��y����O:Z�;#�HԔ=��w�"�;��ex�v�uŨ�.Au5\]�G%�+�QF�åJ))�c�8_�p^a6r�	����#'�Ï$�4���_��|�Jl��,���7�8q¦�C��M��τ� �Fi69�-�9���%z�V`�mǉk���aX`8���Kv��1��[��mp ���n����p���?'c��0g�n���s�����
k�0\��k��@�~������+&M���{7��pǎ�0�x�Ο=)a8��[�&�?�V,����H7c��k��N���4�Y�x��w��!�]��[0,F�hk�ō�$L�4n��f�~�A��0�#���5?�*ږ�-�c�!�ްp���m L���8!���Xw	M������K`��Y	S%� �L�.Y?l1��D<��1,� �v�Wc��$�eX�����Q��k#�;��ь���A����ҍ��F(���D:�������>>��>��:�� d`��n��HXDD]ν��d�_m��0�b�jUZ�*��.��޶T#����&PJ��������?��.�1�{ D�÷��a~2㥅)t��ҧ���U孀�N�f��Q-�q�m�5{�:#���{�@a`.�G^J ��8M����*����F�NR��k��C?�)q4̀���w���*7���k�~��������g�IaD�Lہ!1`�<U_Dr�@ܪ=�7ɔ𚪏��"�^��@�[1T�Ɏ����YA
�;���az��ko/��FBzp㈔E���F��Y��
c �T�HO�s�.��#zU`��V��<?m8���8u��Q)�r�
&l�!ջ4��=/���3�<�ӚF՝q��D��lj����zX������/�[����މ��ȐḸ�~y������A�VT�MȞ�ߒ�}���U_�J�]*qU?���g�J��a�K���=-U�F�;�5�����\���Hɗ��-����ԘíR~u��j�Rc�n�����0�B02��F;�~�2����c�"a��,�#=�*fQ��:Ӣ�D�����S�y~���{���#'|���~S��fZ"5��H��'q�U�?��g��S�(�ך�u�r䙔iʔ�SF���w6Y�}�M8Tt��7�Ӄ�Պ�=7	�G�$	_�L!{�11S�ʲ���$���k4�m!�`[6yͳ��9ݿ,9����>'�\a���sD��Q�y���ճ�p2�e��ֳ �����^m��7�i�/��v�#�XH��)�E�j�u�z��³�@�9䥪0��c�2_�� S	Sx#̓2y""��;.#���]ܱ�;.��`�o����@揢ޥ|�`?1[����=o;
��3V2�Cc(����L�&��@6�6'�=���]Es�;������>+5�5�,D�������1/�v5�t	�&~Tv��E,��Fv�v��X�
K�{����4��e���}h�V}�9O��`U.Ho���B"y�L��O�H���Q�el����к7������sl!�Tü���(2tVta������%�l�E��#D��1N+�\���_���n���U�w��/�LɓcK;pD�j�ē*�}����1�A�ݑ0��VM|Փ��Vn{�w����1���=4,TD��olc���3����n#�Vk޻z���塭�#EP=���7���2�%�w	��T��}�g�6)���b��Z8�{�uN��/�� �����������9J5}�R��x\J�To�6��5���N��l���$�m)��5g;YH��֋)
&�xV�H��	}�����]��%?��
�;@������l<�C�Κtf�J����
�vq��U�Ҫ��}n�����;:?u���5U�5"$+D��g�h+Ґ�ԢD���oV���T:��SW�N�{�ٯ�{Z��.G�UR孥Dߞ�iQ�m!�oa$PJL�w��"��O��C)4D5@P��S�5��y*al��}�fV�)b�St��V5�yC��
ϿTD�}G�>>p;I>ԏ!�5BwX)7�a��W*&/��C�Eü�~B��b�G�`�P�ܑ6�E�m�A�L�R��{)��mс�o�YR��tJ@�z�ch�E�>��BZ��4x���f�x�P�6m��߉�LcX�<��zc��SH����`����P�h��v�f��o�+��hX�wJ���@�m�鑧��^�G@}r�qS	�]MTQ"sŘM�u���y��h^>c����Sκ����և55B�w�Ƴ�����!Rx2��̀��8ل��u�\%?�pO�UL��B��ꯝ�Z�����,��7=Bl�%�i�۸���K�*g�]��*��M��9U���U�����j�ϒ:-}���pr�͠e24��U/Ug\���)_��u�����$R.�s�}�N^�7���Fɋ$�;b��^3Sk���"�F:�_�Y|E�����#�<k�,�M���e�(��:eu'éu�[E����~|���Qa1u�%���Db�������G�]��~b���1��!��x@�L�EM5_��ER=� �,@�1�1���<=j[�������\hw�8�����������%N�lz�{��]2�}����_�EM�r	��R��`�&&!����NE6��4�`YE
�Θ��	~$��H*RO�k,�¾C���R�<̶@y�j��,�(�ҙU���7ݯ`�[_����+����M6<��q�O��3OKUP��M(�w�c��)_�Q���5��Ce���q8&�`���c�h�͸���B�FYym�{�o�b�����ߓ��`�eU^6׍��(���wCrс�&U�ۀ��4Jbl���Eo�QN֜�;��B�إ��}p��}�n�Qm�Ԩ%;^��gȣ��/�|..4��������p����Bn�i3Ɇ>2`꿻��szQ ��	
7S�G�}�'r}��X	��HK޺A�lݓaz�zPH0	���7�	�	wCK�U0,|��7�����V���-Q����U��"�Th�'z���/&l.ν���Q"(��uر�o�ąLXM���n2�>YW����|��<*��6����/�`�������̲]��*ߎ�R ��Sy�ղ���Y"㍩�׷�c?k�soH
~)KFx<e����9c��"�,n�LC��l��qb��#`�m6��`��\�j'�D�.���[��}]Z�*5�K=j}��U �Jj��z{9a<e��}�z$_M��iۚ��V���Uo�ٓ��S���_�f���M�إY����,d�^N�՟��1am���oQ=y"���v���#3x���~5�.���]�cTK��-y;*NU��8"�e+{Y�'������ܻ�����"]�D\�Z �,%6�xe�UN�9c�U���Q<�oN'u���p�S�w������L�'�_��E���5�uݜ�4�4����6���/69Uy�]���{�k^��s���PtJ��X���6���1�MW�XA�K[3 �)����ܬn5�s3k��ZFF��aT���=��<ԍ\�f�۰P�P�/{,xĀEe��=P�Z���8��aA���6�ʸ�NJKb��\�͛���Qu�;����m|�~#�Sk+�G���F��b�h\ūOU;�N�f\�tj�	�=��)~`���y��@Bɰ%� kfr�O�r*�Ҫ�Տn9���\��������]1"DE�(�]���w�PZ@�P��sSח�*��^Lݒ�=Pw�64<D�q��~0�5
~K�4'��?U����ݕ����RR���m��"��pz;��!x�(WEɜt4u2����	�
�{������ZA.������R�uN��M_����!�u���C�k#?V�����ί(�=�MvµބV>~������h�S2oC�U�����/�z��R�m���36��o��#��~�τo��e-gS��;a��O�|n;8�'�*�gN��]�4���qW�zȏ�$�x�QA��rm1>�ZN��xo��V��ΪW�� Z��<J��B�n�#vx!� -q�n3���Lh���[�%�l^�Q<�����O��bӃ����U�d��_,�v6��ittO�l�QM?u^�&�i��dgg�C���E��Mໜ����1� �P����f�-'-�pz<6+y��)��>����1�f��q�$�� ��s���#���e}�S��b������CrG��T�z�{rU8`R����<���.d���֋���W�m�qZ����1�K|D�1���V+j!���E�Ү �ek�O\ʰ1N���S����Q�g�>����]ߓ=��N��]�5��RZ�\��8���}�}����%����&h�{�H.y��M÷����}�3���i��(ǩ�A�E��"x��U��YbdG}AA8�ˊ�Y�=1E�*~z~��Ԙ�	�)6�q�{��%h.�3�A:� �)���VE��(k<r�$L��v|:����u{D;�7�/��Ȫ+��lHeH���n%g�6�$�-�HM#���}(L@�I�?�L,26��cD�'�լ=�2
Y���t�N��=\�:�������Q�ڟni@e�Xv�3����T<=h���~��|�\:gR	W��"w}a�N�~~]14��J��q����5�k8�+�&�4��t	��4��ݟ�6 �;�@V�֪���c	L�ӷ���K� ��d���=$E�����|�x�o1E3�R����,[g�SѶ�|��x�ANYޕ=oI�m����)�,�"�Te� 'oʵ0��>A/{���'QĆN��ڄ&Q6M��,b����^���-�Ejl�;��JtԢ�޼�����F�0ҳ6�����Ƶ���B�p7���N�þ�����e헩��B
l�.^�+y�����K��tXnhR��磻�4�uG�R���qN�R�%-f&�}�S�;�;ya,����s:'���ҩ/H��qa��k1���N�e���a��WY�=C�!�m�����|�$���L�v�b%K'��'q>�������9i��)1g�!b�χg
�;�΋9��{n�I�ۡn�F+Δp_9|cӨ�yc�n*m ��5*��[��?�d�{S��6��>b��c��C?!�xj�U��߽���\�0��I5����P1�P�Rs�����VRHM�u9n�`�#{�q������.�3���@:E�D+S��V[�KA|��(��f��&6��KV?��3.�rm�=��4��܆֣��Ǜ_e�s����;U�k��-n�CPĞd�Iz�۟!Jh)�UO���)'���=^��M�������&J+���CBgdl͍;?��x�N)��Qu'���T���x�c޷�ĂHc���C>T	�>Vh�O��ۥ��m�U2�F3�����Z�$x��1��w�f�c��<�I����Wc+Pγ�ܫWO3�!qd��	]��$uZ��H�CS"n��h�����fz+���@"��]��;�x^�9 �c� N�*M�D���1��6�%D9]�Rc�{��'ʊ0J*h��t��L�?�Gl7�q��U���?�˗RoFQi�ڹ��Y�9��d!�Ĉŋ�a,���`��)�|���QPlv�l?���ޏp��;���Ri�
������T��t�̚�I+e�P�p+p�:�&�����D^������u����˸/jD/,�t>�}L����V7�ղ����5ӳ���Ǥ}\�Xw��$�l�Z��0�y}���}Ƽ���'��F�'���!����"*M�Ost��B�}h�Z��w�?gj9��B����-W���0�U�}_�I�( �{���1mi��a״�S]9Q/�(m�8�N��Q�LDq�(�S��3R����u���ED� ��o�AK���M��5������5��9�|���.t�������~|qہ������]7��,�
�R�_(�sd�I����D9��aBBx�*LR}Go$����:���c�ŀ�Kr�^����NM��&���c!zi��*O��2�� ��1������ÀE���>��Xg�i�ݺ|ao�h�sj$ eO(V�sѓ>%,X��J=��ȧ!�6�1�����>v{�Qtma�����獜�l���J�9}cѯC��1�xf}A�?���r�QT�A�_��>�l�����q��`�O �n��V��H����ک�J,�d�����6�ĭ�A)�ӿ?����]辦4@D�^�MN±y�r� �ϙD��Z���͓w3U�G3P�c��(]�B����4R�<�*�ި1�f2_7���U_ !��Gk͓dí�«3-��^}BXQo�t%-[�Tkimp���n�����EY{� '^�]��G�>H��G0���C�C��#�����C	�J��p�Ѕ���Z_G޸���?�3s���Ң;7�d�Ul��j`!鿚�S��_Wd^o9N���h_*LN,�?�~񿼉��,�y: �q~$e)T!WrQ!��[r��/�sI(%��7���$���.Pߍϒ�ْ�.�m�df��$&�6�:��m	������G!oIE��̎�{�`�ꙕ،(�� �J��s#�|��	�̴?���l�"3J�(��~6!���gl!����E2_�c�RZ3�xyW>�W�9�t�	V�b���;�}Gi[!��3��O�y>�ؒu	#�'�{<�Lm�p{Eo�KM_v� �Sɯ_O�,�S�Ti8{�(nn�>�&���q~i)�|����6�3}un�ЋSt�?/�P\�0���g�Z� �ՏR��#���Bi��e�ލ��u`!M~�$�r n-'\��W�h�烂�|G ��fo�f��ݮ$�ʹ.W�%᳦���!�o5���jci�9baz�����JuEx�7�3J��(ˢ�v�K;�v.Nik����SLߞ>8\:����� 9�g������	NX͂ha��5�>����2ض,9�����aY��z!�`�$��'>?Y���,��8�'U]>�
0p�J��]�o�_�`^������@a0�߿��'��4�΄:�� zG1�������hR���u� � gc;%g��mcĹ�D7�}�j"|r4���8�)���RS]cS`��⌢��:��X��9G����#��?�d���-w�����L��-�
�\���A����|�A<ԯ���5W>�x��1�^������"�m��
�J��ѯYi�_�u��j��8熍���;��F��'N�#���H��攕L�B��� ���C������$\�`�ɘ� �J�39+"�����(W�O%y�j�J��Rw2'�
�p�3�D��>q��(K�	|م�T�ajƕ)4?��fi�S�+p�mm�:c�¦L@F=R>���h���h��%����a��a�YefQN��:F?�Q��pN�'���!�1�n��Q9;�^l��N�)u�i�x����עL5؝Y}�$��V��x���+������,0o0굋G%Y�h�I\��k��ĉ���l&Y|���x�ͅv�
a�u�a����,JCF֙iI����4�	K-C�[��m����lΊ���G�kjc�-�T����GG2Sª���O��Nt����N�
#�V�jD��Y�ڛht��{���S�ud�K���y�|7*"����T4���Vg�mJS�*𨭸H �%)�Z�W���4�,���C���
�.bL��6qMQϰ�moG�H�)9S��D"v�J��%�Q�R�����p�V���#ꦃBu�R��+���aY),c��1����d���D��UN�`��2Q�h��>�BHTFBB���oYG7����C�k�=��v���?�T:ì��@����j��W������-��dE%M|�Zg^	�͜��<4gzq�ZD�n�ԏ��>nK�(z�5�ˣm�-9��\��Z{/�u ���f�01����q�R_�
����&��K&(WR���Z��4漖��q2S�ۺ�\���~�����K#���l|��-E�'�|�!�w�`�K�TU�Y_�?��qfO ���
s��ӈ�(��$Heܦ����h�^�.�C.e;.���	�b��L�L��m�sA!#��Y�Н����j�c�I]:���:�Ȗ��������o���)6?���A�$zҐ�h�qÔ�5�}4��������)=��Ue�/n'������-��xޝp�����L���BР!��57u�b80���@#���ؗ���0)�r��Ak�»l\E��⑻w⽛)��HP�}���$��NH���`PT#Za�VT�~)y�̩X)����d&�J$�MH��N��<�W8�s��h57%��d����`��A1�՜~��>e���[ˏ�}#{M�[�'ż/3���{~�y�I�������b����"-���nG��!���TG:�\(��d����/4P��Gj�5�sXr�Z�"�Zж�X�\-�Xc,p!�/��A�r7�����e���֒���	��1����Zi}�������0�>AX��ڦ�χzja��8nXҶKr^R�B��#)�h�`�Ҽo/���wTr�4\�D쏣D~��q�8�H�}Ҟ����X+��h�Ԁ�b܆��>�2/� ����J��;[uQp���z2���6�j$Eal`xzV��}pA�I��KI/ 3�I��T=%X���"���W���c�d��	8�R�~B�)���<��a����@R������m ��o����U� ��^�%�_	q���������"بQ���ΒL���\�P�X9	rJA��"� ����w��X}�J�@>���4�=�/K��o��U%z
�Fل�7|�
�����d��-�����0}�d��4���#g`Q9�T��䡮���xϠv��!�R矉^��S��
W���cX�Vy!)���Ě"�iI"��=�Yڇ�e�h?ql�Ji�7%��.v�"���%�H�o��k@�S�V1������� v�	E��̪D�Ů�k�_�U�dv�TZ��}��n��ʢ[_-��a-������'�>y�0<��,�����\n�19=�_���u�1j�I�@����<N%ϵ�'�Oat$j��R3	������>�M�4���\U/�t���O��ϥOb_,�Z$�r�q�;P����ҵ�A\�u���r%��P���<�g���ކyӪ΁��4��%;���5bM��ߑ��e��cXԫ@9�@�ԥP��
�ك�r�s��'A�Ӣ�[ӝo�_>�>��7���-�� Y�	�pvC��Dl�tw}e��Exat��2��x�4z�M�;���w�㽨71*'eeqI;��|*�w�׳\�������|>G@_mY���-��L;9'�_<��1�>�8);D����.�
�b_�V��p��R��t�f��*�Z��PkA�^tS��}�nt8_=�
1|y�z�ΆgV̈́q�����p�tCx#�FreP��a⬽�M�����Y>"�a��@���"�>"������.����[��j���!�T�n}�]�"�k}T)���H0m����������x��Г�p�	��S�|�r5\�	֕m��©�5Ro�g��г�5�C79n���T�@����C�o$��u�����0������ݹ?w!��6,DՁ���WW)��}.-t��p/��{/�����"qo��1��
;�M2��C�s��ӣJ��T�q��yd{�-Bڛ�������R_T��>֎nH6I����6�A�~�������hO�5:�	�vy��9!��a�@�C6����Ɔ7�o�뽕�-�$��v�,��Ͽ��&��bDTB���a�5��$�.���ʭ]^W�[�S�uy?<�J���'��~�ϙ�m�ί�>���u�7#���W����x$Ł��C�,מ���i^E ���w[Ԧ�ͥ�3��{x�mGo/m��cE��1�C��b��b �$Ut�1�����Qp�{�Z�������g�yH�D��=�\�x���{��m>��C�2���iyl�����\1psW�Ӑ��#�X[1w�w��u��&��f!֍�zxDjIv��f��40QO!�$
�CopJA�KK�b�g�����|a��*�'�&��S���;nW�w�&_��C�kW]>�}��.�Pu5�u�6g�Y���M51r��ջ��jڅ�����hn�Ch��WI�P!-�3�p�ZN벅�^G�j�$�D3��og3�U���7�h���dE�������+Vw�?,kFF�mt?���+���yrfq�p�R򲀧x&�.�(F>7R4[S��jA$�>�5.1�ѱ%�%[_�à��G�Q� jG�����������4��d��εL2�����&����xI�ƺ���$�}��8�Ǵ2�k1Y�S�ݽh~�aN�B��_]:��Ս��ǻ���s^1��~���E~���$�j4�=qVzy�d^w�F��@k5��{*������m���W�ͪv,QE7V�j��//M�Ը���?��+kKWA���)n��'�̃G�.�h����>�bB�{���ЪOX�1���0ܪRm@c�I�O��@�|���*�U�!"(�$�˲��ڲ�lRI��tlY�'�@��w9��|�O����>�x�������o����rm�D�� ;�s|�b�L�Օ��?NI�
w~.�t���{B����;��ֲ��8�{2��r�K�V��.�V��.����c�	��;h�Dқpج���/�Et�yt��z�üa���+�|�K3���x������6�o�a�{�Gn��)�����|�Ei���`�J8?��6�0��pV#�ŀ���X��ڼ���aZn�v��Oݕ����I"�Ʃ���=n�ydb�PЁ�	�GF8Q����X�A2�����'_��?F2{v�C#���N1��&U�8ߜ��Ɩ�kw�cnbl���c���0�`=C�I��s�E��b3"r,o�������Ø�8%6:��W��ki��Ygy����8�?�������Y��e(̞lN5�Yhx��=_"�����bFM@tJE ��"2*�G?�����i�^�Qx�G9J����d��oWq�e���v��7#�y
�]Jĉ�O��9L���� ��b�N��#��� ����޳���r�^�a���z��{	��[���O�r����@�������S	�ҔЎ�8��z�(w�P��h7�㠏��
�����AE��W�U5��a)���ˑ��hv�%��!;�=Q��fO��5���������vS�N>��ո~'2�:t�1(�Kך(f��x �A���"�w�6�G^�����Ҵ۾Z�����R��/9����u�e�me=��3�Ux��R�A��6~ߣ��긖~8ebֿ,H�L�̎��aY������^[Ù���w��0�7����a1���#�9�9N���7HD�.s��V�z"umz�z�VK%���Q�%[�l��r��q������-�ʄ$�TD�!9���8�ܰ-�L�\M`5�}.~|��1�:zS�!q��{�����j7�S���Wh�Myo���j�_K+ß"}��n������Of;��tSf槑s-�x;8!^M�%{���N~A�A��m#`���> �����w���jW��p��0Q3Y�}�_�%�ٕ(���ؕx��i�X*(�����N~*[��H\�Y�qʓ%r�V3�J~���nO\�pe6��ҙ�t���S�y����F�qה�0F�����b~(��:�i:}DvI�)��hw�����W lD�Qq=�~4֠[�\��K5k������c�m1��C��D��O]�Euc�����i�yp�Da��P/4��sxH}���0ž�O9^CE��7母
" �t�W8���H��dk� ��C[�w���7tLJ-T��1]����b��d�t�7$P�b�8]^
��Y����L�	�ц3GRqe���-%��.�ʌ�#>����M�Q]�R1������-
�,�uSFq�V4.z�=r����51����Lnm�qnEw�p|l��`,�HʃB3�1=~$gc��Re�&�A��:�Vfo��5{��`�CB�y"q�xy�,ݛ7�|�B�p�U���>N#�!���)�4��k�(<&]�1�[9����u������:jN��Y_,�s�-������:k���kٸb9�^��y��E���j�L�� 4��k���9Σ��rl��8W�)�5Il��\ѷ ^7�:��!,�,�4�T����j��jJ��^��
*��5�e�	��QL��ש�4<~ �
���38��>�-u��v�{�{Tyt��.i!�����m�]�/!Ӄ۟-��*��eO�V�� "=���z��Tޠ�]�d��u��'4�������`j����8��99�<Ig/���7�A�6����m_�ʖ|nj���Qp�䢸f)���τS��`���N/=�ӓ�rXӘ��2����͢eY��ﮯ�Yu�%�!i���(�9]�EC"��oB��]_��z�����H��`��uq	�4<*�6���1��7���/k���b-a��	`�q�;��hS��]׳� c�9O%��I7�:^c�#7�..ڕ����wĚ��H�ߢʿk� ���u��s�y�4��hRW5�����QJ#�Sb5��Tk{DȒ}��3�R�G�f��-> �@����6�E���'��-�S��4t�w;n,�ٞ�OQ".���s&�]��^��of5��ՠ�ל���r�؆���D/�B��/*5hZ<!�|Ƶfֵ�J�����d�'�����C�;��8K�_5z�G��
��i�l8� C���A�0���B*0�z����3�x�5R�����1��0�}ۇ!BV����U��D�{Ht4���$z4)�S�V����a������G�w�ň0&��WK����~)���N�X��d��U�2��ZP/����'�6�fs&�mC�r���T��?�A_����Tƾ�C��Ǭ"PW�Z丑�H�F��V����CA�q��/�����]M7K�(�څ�y��U�R�.�\�������Ŵ��u����:�,�bO��EL�Ć;
����IǙ��Z�Ijڕ2����t�5>z�GSO�e�w����O�O҆�	�Rgɹ��ާ��&�D��.3Yj/�$��]ȫ8�>���.��q�j��:����m�ph��@l|b�|j9t�1t57H��!�Xa(����/�^�BV��}��E�q�N{�c�I/�/��Y��+���&�(��Ʊ�Wh�cLobW�
��C�le���g�8�,.�K���G�O��8w�3qK�X_Ķ��A��%���H��k=o!�Ss��3�\2DD�7���eM@/�
�	'Fc±[>�-$uYFop��H���5�l|-�����6�4a6�v@Т,^����DkH�������G̃��j�:!u���� =4r����ވ=:���Q<f(��T���fD����;��yRUf�@�/��{s�����f_� >��~Q�ۻ�->+��u6,� �=kk�Υ݅*�HE�i��$F"�u�I�xz��ښ+�E�$D�oCig^�X�L`�^�z�	H�3q�"/
�����|r�)-	c~�o6����oȢ�F�e�.�'tz�bw�K��.�o�C�>����0�_wp�p=2k��!�}Q��� �>*�ִb�%a����f2x��sĒ���w��u�kF���}N4��9�s,�UQ����>N?�rX�%ɁbH�&i��Z�7��^T�Ѹ���]k^�C�2Wڟ������#𼐋 z�)O`��e�f�:�"�O
��"¥�E��dSR(��xe!�l����	�S�jbG-�����p$9��V��]ẋ�,�:	�/?����౓PbrU�T��5q�K>���~����Gsc-���Sr��L�,[l��dMZ�Ql���7�U�&؂��7 �{�0����,�z���OO�1�1�Tk�:�nX��"��T+I?^!t'�86�e���1+V����'���g��E/�H/�c&�s��H�RA�~���h�A�!�]�p𷝧�Ȓ3�����ں��(0 ����C����36�J�0�t�E�J���� E����A��Pg0����'�5��Ƒ9a���;Az{�=pb�27 �;D��9�����0�]��m�y���|Q�� ������CuB+�{1uҧ�R���|��^�tUքD��¯z	fe������$w��yI��WlGu��OPŦ���Jl����5iHM��M|J9)��QJ+K���ֳ2+�%;T����j����6�7.'����?���}�OL��� XW��j[���9$7��G�D�/D�����1d�Đ�|�����Ԩ��Ϊ*��|x�WWBG�0^[�ꅁ'_(ekl��jQ�D\CMC��I�W�5O27��1�@�J+��/|� R��J:�jrJ~ҍ��׊
�B�*�	%��8�S��э���Q�g�������Z�,|���!�yvӦ��b���p5C<o�v��$u"ƪ�V�����%��H� D�_@�
��I����8��xYd���M(�&��
#ʺin!�t9�>O���-��SG����$火Ɠi��Bv�&���n���q��}���"Շ3�zK�U�+����yY֖�x�B��q�E������\�D��ڰ��nǃ�,�^�i�*�'�?�)����C�}=�\L��n�X��|��4 �6�p����6R�I��l���xA�����|C����
�a�.7Gc�v[h�״�#�gY�K)絶 V������x��V�Z��.�n�>V8�$F)@��p$�M
��.$���@A�(�I��˪�;�bK�8�pn��qy�#N����:�J�b2�^I���0�q��g�i�MUZ&�Ŀ����fp?{���0�~����� ʏ
��/	�\Z�a��]���/U|~H��p��X<�H��0�k+�o���xʋ�O	��M}���R�j|>J��u��1K��qY��W!��/b�^t��Fi��&͘=�|�Гh?����=��7����*��cΪ\i���O�o?g&����4K�YJ�ͅ��b&���؛I�?B�ȷ�e�Q�I��P$�{��d-��B_R�&i�h���g�+��]���WoA�Ι>��L�Ts�9�|��Y�4�+I!{pl�Ϊ[p�+��A���Z�cVR��;\����C��Ɨ.����%;ƞK��aG�:&���ɮp�~�r�_H�H9\{������ �-���)�Ћ�����1Qv��l��pD���CX�q&�΀ ��g��r�2RD�y�������0"@˚��F�v|Ȑ�9��]�����I��럲���A;��w�3�zD�Ǧ���q>���,.�E�;��vf�Y�~e_x��<Z�g]V)O��N�7����u����¼%�o��K~ː=�wV�OC.6xl�����;HB"���5��g�?C{'�i��jE�:�>]�R�I}�K+:sV�$ �N�2 ~�d~&�څ��C�����/�	?�2��"�bF_�e�����pF��ΑP�ǿ���B�=ܯ�q���U����8���D��o�c2��v_�c���D�"�+F����!/��A���'?�蠦��0.یOށ�~�P:�$N"/�5��Q�=�H>��yD�X�?���y�QߏAi�f[[[q��9���tz9Z���ܷ䄐�
&��'/����&�8:uKk�Xl�������L���,�h>V�q���{��DJfܟ�톧2���/G9�R�0���Az���V�c�6*z
&+>"��%�C���������[a{�<}C��JF��-����k�����-�h��t��'���H9ԛ��8\z:	0��Ӝ��8b#�����
?��Ԑ$��P���_��aB`)o%��ѧ;�g+���T)�R���>�������/j�/w����19Aې��^���g�w�����D�I�uO���v��X���(���G�R�1�ax�����KZV�og/�!�؍l����ǱG-�Ҿ�s���2�C�^~�	vW��G�Gd��}a��d�_�8Zj�UA��o$
���G�i�Ne��c8�T�=�<"��	o��\7�k�ʬ�J�m�ɵ��`�������[a���ɟy}��Rb��i�Iz�����|y��A��(sg�n�5��sF.@��@�m�ԃ����UL���8�	B�x5��&y���w�~�pߝӜ��t�߰���|��(���r�_�Y
>�2v#��]m��r`����{=�y�#�!����V	�����% l�A��~ok�r�n10!���d�(��]h6����?��|��q��5�c������vQ��{����!���V��o�?��D�ykR�$qeN�h�p:4�S���н�	�@CW��PP+����^����j���v�� ��P�]��������_u��3�͋Pb��Z�抇�T�Ř���)�+p5���<@ÿ7����`ټ�X�h�,���K�����ؾa!� �~��_�,Ɓ=kX����]�{����*l��3vlތ��f���)Ե�a릭D$1�stl�2̞��E�ǈVae+E� 1S`Oq?kV�zXG���(���>v�����!0<	����6*V���P|�@�V�T'b��LZ�a�xiZ�n�	�Pq����1�˰P|;��F�b�nj1��[��G�+h(����KHt9/�(�QL��O�@i�	>c��E)�/yU�7Иw-E�А��Zb���y<<ŜD��cȾsY��6�A�U>KF���}v�Q\�)�.#n�t�
[C���,��>���aG��\&���x��|â+��1,��H�
�J�E���b��*"���&$KM��
KQ@�+������|N�#�'L���#0=.)ɗPW����|��e��5��~����DS�*��ó�xz3Nmã���sTW棸4�E�(�0\D����U�\���y�(��Bn�+d�x�/�����2���u�R�d]%�4�x��!F�=sx���{�d�Yc��B`�f�M���-ŝ�a��_)��:���Qư�.����؞��V�31ؖv��k�D	��b��~���i�����=v�0�m�=6�g����[�m@Z��;'&�8����"��y�߳��6���O�T����h�~�����m!��?�x���0�7�+n�F�"_{���n��DڝL�2.�ְ23�=�oW8ٙ�{���wbݚ٘>u1<�MÞ��q��!x{�`Р!�qp���t�aSb�#b!"�C�|�2,�?"_İ<&�D�S4ç�JZ
����5�	u�hk��{b���df����⁘�)<��Ǧl@+!��P�}W+���*�����;���B4������ol@u]-�[ZQ�؂��ob+/�P�¶�M+긭Z��&~'���X�|%!���H\�ybH�7o;X�V���M���0�5m���:,ں�a�
���!�%����n�!����#0�1Dd�*G�������X��aY˰r��!���栿�Dt3��y����e�:��P71r�l��ρ��4�!�{���r�!�A�ȭ���"�hV`�+$���v͗�c~7��lS�\��\*&��M��%��p}M�P�r1!aX�����2w^fg"��]�8yA_�kV�Ƌ'�PF�e��8�6xM7�@y�T�@]�S�?`Ҙ;h�|���Gh�z���h�~����<�	��C[:�j�����^���9*��|��{/ԇZ���6n؈��Bl߱��6���)�)�C�Y�C��Ĵ�b�잖#Ѓ���0��dїX�fԝ'�y,��Z��َE7c1\����7�:�<�g�	b5��R���Į���m6���F?Ǚ��`�4�=���e��!�5` ,X��ش�//���:�^�D�{�%�{Q��هP�|2����7w#��Q�?8�ҧ	(yJ�>:�g��GP��(J�c����sY��$�����hz�͹�xx�:��M�p+s�f�V�<~|Y�$����F��c4~p�����Fk
O������.״u��id:�+7m�m�\�d�N9�OJS��R��_Űxn����p	�c�0�5�11Ӱa�Nd�@�4í��_W?���W ����x|�.�݆�K����
_��$�{�<&����(��!����B!,������X�G��e��w�����-��o����X�ʲ|>r�~0sp�׈q���~>���m�
8�[�O� �,���r�v��Q�W�X�W���ZD+���b�5E:1,_G����G���	�b�
��1��	�v�V�m�J؄�0l���p�"����g��*Ɠ'/Q��V`��T�Ǆc��8��Xc���/0L�=uD����������j�y���Jw���C�5��>/)�EKd5������a���������]�a��>/ǰ�:����0oV<ܝm�~â���Ɇ(6F�8{Z\@73����S�s�z�9qgX �3�ڃ`am+Go5u���(xG-A�ͰZs"�$b�1��߃a��BJ(�K��"b�eY�	_ӰEж�Bh�J��v�@e��/3���UhijE[�;�U�◽��GgWlݾ��Eh���"&���"�������]������5u,]Q��P��]�~	)�Ҍt���`YZ.�jiF}S���p��E"86��X��Fd��/��n ��	��Vb��u-�&�s�:�j�Y�FN�>�Fς^�\f!!,0�����E+���)����H&~�h��� � ��XM9��e#D|Į����aX
!��X>����"�%����s�+�����)km��R˰i�����P�C�!�/�w��q��V��0Al%��@�� 1l-����Z�nE�H�".�S�r~�RK��9��.��K~[z^�Rd[�g�nK���ɑ,Z�Ed����(�8-1��Z��4{^d����Gpu�����8�w��,��Q^����,�Q�
m���Z��U��XqՅ��X~-U���#M�\�'f�KFE~��/���!}��HEI�-e�!��K3�m۱�,ѫ�֮Z���<l۶[j�o�O�|��,�]�G@�"�-���a�f��"?����F���p���Sa������E���t}�4�`��4�xO���l"g��u&1<�(��~�s��j
��p|?�=��C��
���譥'W+lڸ/�&���>jJn�g�(I?��"11���?��;����J���Q� ~v�9���'QD��<=���'��YTe�G!�y��'�4���i�W0o��8Be��L��{���C?s�A$1<?8���aq�a<cc����'O�bB"�*+�~����h�׶	��F\E�	��6�f��+5�2�{�rąx"��b�i�
�2����zn���	�����+:>�������?6n_FU{.��	ߖ�<�<Gs�#�����l�����	$'����3�z~U��!�+
sP�O3Ź��p�.ә�(�z���'�p^?KC6k�|��ª��(A[S!a,�	�ٳ�������L�<֎���s����3~<�Й���ep�����)��v��v��c���_�h�%��D�a�v:���(�+l'0�5��q?�~��E-�Ao:���S8��5v��y���_e�d�ʊ���&�G`�ܩpw�ò��v7U��ȩ���C�o]O�����%������Bo� lX�
Ey�hm��~'�Z��V%���~�/��t����_a��j�g��b��pq�&��Â�"7'[�X�c|t0N�܉�ۖb�Xlf�y`��8z {v�D� �54�gh*�3u���(���0a1�X°)!,��U�o�@���؈�3	^��PY���)�8�i�,µ��k�X�բ������,ӚZߢ��n���3ahf���P\�����/1AG�l
��r�eH#�ϟ?�¢l��8��gY�ȂX V�<3�7o��$	���QZY���Z��U��ֽ�������1�F���[7������++���Y�V5�����S���w��?��}��*�:�Y]bX�F'�
K�������WD�^Ee�J��,�O�~)
��0*&�P��*0+!W���uŌp���5����QL���n�&��Z����<"��]&K�$D˰�a��a����[�a>30�k�4;]wя3�̂��@��
$����2�-��e-��b�7�®�C����TZ%�~�o�Uw�b=y:�+�؞!#�Hh�H(V�X쏏�p,��X�~á������G/��֝{pq􀑞�A�����
r��(�
J󮠶�*膢k҅aՅ�(˹���Q]��ƒ�溅�N�<��Dr�D������4F*
2RQS�U�ϱy�f��@OM,[����غu�AE°ܙ�"�!����C����^�����LC%�:M��k���S��~�W`���A��#Y9�� o��$��}D_a��Pq��^.s��y��8��&���z��k��z�P��E�Z0�6ǂ�sp��E�g=@qVJ2n���u�d�A��kȻ��̻���v��O��`.{u�9�bb7��	Y�\�c�<�2b�$�,2��ۇ��wyi8s� �N����t]1��<g�[zC�!Zn���~Q҅�?�2�ݝ��I�p81�-��ĉ���xURW1���8+w�̬��r+�RH�Oҡ<Y���a٤2��Q#�ܸ�9e7���`�d�i���<�L"�g�w�L��Ƭ�K��!*3Qߔ��Q	�.o���:��]�K�W<B&ko�ǓۗP���T��
)� �3x��&�_�0��y�/�	1� /� �u!�u�<A5�d_����5�_���"4�V�������g l\�a���)1u�^�_��3D�up��aq]W�*Zi?A�'��⹯�s�|�a%xw������;b�v�r8$�!,��aCb��7Z°��$&��w�%�Ux��-�;]�!36��M������{w�#�܉�$��A�pI�gq=9G��Bx�z~������ưA�v�2�dr�����A,Z�ۛ����ĿZ�{����F�B~[�pc��1n�œ{�`���>�ΰ�����H?�?����K&a�����.>�K�-HS����AC��:;����1>�� ��;��Ba����l��z��/a؀�U�P�a��E0��s�	ذ;%u@M�[�WV���5�,X�������U58|�<��ada�����N�]TVW��kBK��_�*B���n���(`�����c���Q�aV���.'�B��;�5�J�#J<|�k6l���=�,-�q�v�TW��m�E_����,!����P�؁����'�C�b$���	�����������/�c�����_�I>E/q�7a�S|v"TB���u]W���� V���ߔ.����RGkz��r.��y�p�"]��i9��0����Ab��h�E�H�@`���TD˰%1,E\ B8��a_�4���@�@���q+�.+�T0����6�~���|^�h)Ҷ�V���|��.-�b�H��d,��G-_h;�˓��1���>nܺ'bX_����g($��ň�I�+MEc�-�^Ce�e������o�Წ(�I@��p�E��
!|兩(Q`��.z&aXc�%z��d��9زm�KV5�eE(H����3"
+� qA&�����0b8�,#��>	C�f`��T��x�k?���[}�a/|?��#X!��b�e�ܦ����v%~�硧�<�x�8�E?��P�1���+T���G�������d������$��<Am�s��&��� ��%d�?���c�!v_�Fi�y�e^@�˳�c��H�}r�ϋﮠ�5�<������M�p�&�B��:h�F^��Ō�^�MV���.#��ơ��@��A�K-������͇I�,0\.0܈�ʪ�
bE7
�-Tj� ���`X4Q�����r�]����:i.'·KD,<�°��/(�N�I"͍�R��MO�^��y�����ԾBY��HK���)(�x����(�{N���yJ�>fI#O䤧!;�����e<xk*^���'��|����%m�E�xSAWI3:=��cFO���+�|F��5c���YO j�N��o1��|���_ﯥ+��{�-��N����1D�@G����0���3g�����E�hnm��C�0x�6"G�J-���r���".�;~x��׮`��M��rG���������8�7*ˋ�.@�� -�v�����_NW���(oG\<�	����0�h-])F�ps��0<.:���?
�b��uH8�N��5+0|���f'��l}�k���:y#\F��Ed�[������
��qsb�i$��0���QVjZ>H]�X�5�,Ϫ�[!�le9�*� ���G8��a����t5	�E��b
�j"�Μ?���\��5U�k���e�QjV`���-�pCk�4���篱b�z�����ѱ����K�}x'�+�n�AiU*�P�ЊRVZ���'%�X��,a6��Ӥa��!��_d�>ǰrl��[���
��Zİ��h�	�'��$kXF��AZD�i�âex��lh8LBӑ��(���-�#�p?��U0aJ��0l;Z� �'X��Bx
d~�a�S�R��Bgd#[H3�Y���:w��R�?KW+CX
�/��P1'*���'���܏Z>h�}#D�O��W�p��]8ÆJ�'����b���/������ɿ��lb87�Y����]2K�~I�q9D0!\�e��3]Q$�p>1\]�U�O�y�&b�B�&�t�Ûb+a��5�E:+E�t��Ӗb�1Ӌ��b.����Q���A���3���������aOb��v#`��>S�X��OG_����6=�磻�|� �Eq���<�v���YY3�D?#'�bF�ՁP�Cc#�L������a*�r�2'���[(JOF��(���K�.��#��I�?:��g�P�}^S$Z��rq/�%�2sKVχ��4��pC0v'���n�~�~��J�(�u�Hh�M$���{�	��1���{�dl:xX���;��aɮL'�� �W���#���:�x�{0,=&�O����o*�U�����*,Y��31m1FL[��3��Qq�p��)������~CZj�����w���:�Ӂ�|�#bk�_�8�!w�h���	�s�0�!|�NC^�]����{(+|�Zn��&�u�hn�FkAܒK�¢5Z\,�@4g������q��S���p�Ô��1e�1�؆�ٻ�9e�R	9����%L�W�Ls"R���pg��K�1���FL�Yb8=� ����q��~��BH�/�N� /OG,\0O�E���s�.]8��GH�&�]N����ؾq}=�_�'z|�ƌ���O��o�J �4�Kc��i��z!�<�g�����E���$�n��3_=ƲEs��`s=����!쬍0)&	��_�a���޵W.�1�+Pn.�PSW�]�X����K�&������>b�'����×��|���İ�/�wv�Y�(��e"�����d�������ߡ�}�	�"�iEU5�jjCmKҞ�Ƃ�a��GOoL�5'����J1�Û6�}���!�(M<�k��F��,t�Yಐ'�w�����V�� ��M�Z�.�^04����p%������n����ʛZ�
��ʑ�����A�����g�'u�P X�eR��|�X���C�����r	��a+��J��~���l���eYB��0����]/>n_�Mb ?��h�$�@�==�a5��� -�p��#a��L�v�L0G���|�]s��E��"8����e���Ī|$�/E��D<	����@�4�1#V@���մ����()����(��ğCX�?�ڏp�OZ���t�-V>�{���Z����.��SD�M1A��y4E˰�#��M0a�<�x����҄��mGe�K�U<!������kh(������$�+���+Ҳ��y�&��<5\��"r�EIv"*��)��	�y�)�*zD$?¦M?K��o V�\�����{�L�2ؖ��B˰`�|�aY�����X��0Jj�5���~3��8�u�u������ý����}��YA����$hx|�p�y�F��&�s�S�.���N�P����1C��X��犁&n�n�!,�u`g��S�����r�(��K�>��Ҽ4Ԗ?Fk�K4�>Cu�}T�=�����>���RE"��U<����'~����aff�AK�t��m���U 4���౥�Ϭ�U���h�r�Ji,1<��ww��g�����g/�;�K,�ˋ��L��TV�V��J�Rj!��#��ƕ��1�E� ��G0����"�s�c}/:޽C~I9�o،�fa�Tbx�rN����S���YS���m����R�ih�y
��KWu��=��x��b�� �BC9�[����W�)}���g�ST?��U�O�X��_P���&�UL�ܚK�1�<�Z�{D.؇����v���hxOGD�ĭ9�1��7n+g�[�h&J�F���X��� ��8�������*���(��bXt������#�p��y<�����y�gx�Ё��sCh�lmL0}Z,A���V�KNKI]'Μ@r�y\O���[7������	7g<|po	_1�֛�fVL�$���1��a���tK>ߖ�eX	�Y�O�d�,�XK1��!�Z0�ӑ0|1� �˗M����p��Yܿ��G����{�`��1�����$�|&�#b�G��M��O0���a�@	�b�|�+��aq�<�u�:���7���1j���y�y�9��K7n!��}T46�����Uu�iy��o�|�f-]	��;�aTl6�=��� ��w�>��˗�]T�F�5����f�qCSRo�F��T�@�q��S�=pS�̈́��l�O��{������ՠ����߈��Z\����G��m9�g�M\��i��}����
 ]��D�����^ޙᡫ��Zj	�%�����d�s�%.*���A��\�(V�� ����|�}�\�y�?��_D|ģ;1�j=h���n�|XF�<���΅�Sz�������AŌ�!�İP�r�ل�#�>�`+�W�"�i~�j���Uъ�W\�/@,ǰ�m�`M;V�a���۔-����=,��6��6��ry+��5�?��,�;-�~G� �7�BC;��#f�l<�z�[w����SCCbxJ�H(+�K�fK�!4��F]�MT�$���ȹ�r.˳�<�P�*�G�����(�NDqV��ϸ�ۨ,�������}��?���?A���_k׬GEE9	]3�l�������%�˺L����@�J�1<��/��&�{����z��p��&İ�o4]'K�(c�{�[����}��N�.���0��u�	��@���j�S��Bu�)���A:�0�7��h����+a��q��6�;�׮���;	�u�<n\?��`�n�|̞��Q��w��Ơ�親ukh���������%��d�]b1�3��S��{�{Š��hf��v,�l;=$O�o3����_p��Q��,J
��>��娭� �E��,��g!�%ϵr���>�Ҩ
K!xe/�53K ��֊q�[�]P��k~B�9�� �S#$n1FM_ �Q���֯�s��]K9j�چ�x��oEҙL�o$������0n)ć��o&l��ސ���L��5�k_����4f�ms&ڸ�n����[���í�fI�3�<��##`��7� x�� r�:�/?��ٻ6k�����p�#B�1<A��ʆX�>tBX,��� `�t��o��k��2���N<��������6�W0��[�ѣt��5�-+3{���`-88YI#I�B�1c��I���R��y�;uW.�����xgŨ����Tܸ���q���/�	wG��em�^��*�]�&��a���K��-�Ҷ3�)�I���N���l͍`0l���!�p�/;V�xY�ukg`�/�p��^����}{�hO���0l��=/X�E�=|��W�y�
X�1�Ɉ�ݘu�!�mF,�E�TXL$��4>�g��ᳬf�J �hlCqmʉ���\��6�o�(8� 0j��-��]{�~�v�:rYE�hhoC�[� @�2��^�.q��ݼu'v�9��ֱ:N�����K�z�ԟ���� nE˻UW���[�y�>���n�q0���)�M�ϗF�}���.�����^�*�X��:��b2m����t�Dqg~�PU Xi�ke��aX�����31�I�_���b�xt3%��0Wz~R�-�e��E0Éf-1��E4z(�}�B�`B��
��aKK�z�N������1�$!R7��ӟ�ˈ�r�Z��{��@'Z9�Fz���Vj)�1c_3��İ��ԍ�id�)�U~�>x���px����R˰�����ũr�@91\�Ig	_��8�
jąu��	�������ř��.��*�����y%�M��i���lA jc���(����u��a���b�	�>�a8T�lb�o<�C�gH-ßb؛�c��.�U`����m�+0L�1��g����r��i�k?�vq���B��.�n�T��~��0p�+wD5C�6���00�������a���
�'��|���G�Y����Ct�1`�hh����z4B_}'�6�DC|�ߕ��Xh�M��J�𜊾�`�ݽ��#����u�l��n��u7{���nb�H'�[>�p%�n©t�4҄�a�K��L'���eCS�,���~�5�Uh��yB��rFM���I��?i§��Ig:BF�"(|$1�tf?GGS1Zk��\�J��5-կ�^�����o���}S�5f����S�_1|Jk�s�~�7M����o���7��h�"~_���O��pkwNΟڇ��������3�2�Ŝ��p�^������c7�b���r�
�*��
��J-�&_�oŰ<��G<����#��C��0<�3��8~څ;w����>`˶M��
#����u���.&N-�&��*�p����_I<#��x���2|=�V.]�~*�����ix#�7ף�n"���-���=�Ҷ:1,�uf^��3��'KS���:Z���c���H�r�ɇq��.�:�{vmBҥD<�;�퀾�1҅��3�B`�(f;���qk��c���aFa�/aX9Q�a9r�ƭ�����s<�>ց��9�����hN_����z�6u��(ilAVy��`Ǒ�7>~�r��Gp(��~BfQ1޼AMs�4�Fu�O¸��	��ab�����?H:��FDb�/����k4u�E_[�Ђ��7h������2C�<��SaLN����0��Z��e?�п�a�k���X~İ�lB�
D���VHK�y��6�0r-,�m�i��Џ\Ct
4.�@E��oİ�:��ʐ��^ß��OŰ�|~��rO�&Ěy8�����p�<Ë�0�D� ��O�&��8��	5����aY7	�E�$f� V���"�+���鿶����R\FB�Ċ�a�b��{��Z�4������hʣn?j�c��1U�QR�f�s�:�Sw�hh�������M.�k�}$هB����6��t	2J�p��S�����{3���@��e�(�"jKn��_�"`\�y��MB	��u����|�J|��H�vb�8�:�_����1��ê:X��G�VT�1����e8*<n�E�B�a�%���`�i�G��߉a�M�T�/���{����w�`x6~p���Ĳ�,���������Q������u�y�:���={fI"gP�9�s � 		B"gp�9���9bL06���r�B_����%����=���٬u�ꮮ���nU���q	��R�N
y#���Lc0�,��	�d�̵��L�&�	�3L��θ0N�<�&�m1a�-�ϰ�s'L7w�L�f��,/̲	�T�`L��x~ީ�y��%j���᫸ߥ�T��.����C�ef���B���|��\�0약;�~f8�	[cK�	ê���m�`Xpn�RL�@̅U�
����c����1܄.^ ��9�0����%��l=Q���K�B'g-Bph$!�]�7�����!.�jo��ՠ��q{�b����v�V��%H>�~b����|�ӣ�z���Z�Y�,C=_�崞�jč�v4�U����A����GxH�b����+ò�� uų�ځ�E#��1��z�t���ܡ�>v��JԼ��Reէ�p�E�h���5�����܄`-�%�:�}�V��/v~)�k5��T$�/�ڵ����Å�5���?�)�L��l�Դ8�����%G��ǾǾo��w���/?������%���LM8��3G�ǳO>
K�و$�����^�LF:�D_w�%�J��b�+<�7�I�o�h��ol�
%#<Z����[����̅?b�
{��|�$�F�/>C]m._>���������*TU����q�7�-��hl��O�O�����'��@x�j$,؆�mpK�Zm$����0c������C ǚ(4��0���v��{�ߪW�xe���Zx���_�*x$,�}h�
�����tS7�����{����v����>Ǫ����`����r�V���A��U��H�h��D'O��(��/� =#!a�������x�^����u�}?��e�O;o m�[_AJ�F���B�.I�T��Cr9?k9��y�R7�2���M�c.��#0lO+���D��)��\� {-z�+^D������cb�>X�s�SBxÆ*
��h$��W=z}���6W#�"C���h�`,��JH��d��0�"���"�=q%1�V�專�1��qi꿚'�S�y�wM�47Ɲ&@��0U_��I��"��ʀ�$K��\�<��Ǽ��㗫2ן	ʜ����l�.�,�6����'b�d1:�ۜ���-���sb����"�*���` 	)�i�!aK`�D,ż��*s�F$�s���+PS�7/��G.�Y�R-|n)Y�<r��c)ud�J`������,�����g�g�~d��bU�
�?}]���V/��g>@{�^t5�W�����EkqK(7��:����a���}����43�>A�5U}���=h�����g�~���}x���a���3̰e���7��W^���&�za��t�F�e�QL�aQ�k������x�x�M�M����<�қ1�aX�P��$�R�W��"�����UDe9�V�ë�bB8h�	(�X��_&����g���a6��P�)�1�-c��p�Y8ƙGb�i&�E`�E&�}�X�b�uC0[�Z&�� L��v�L,&��rsI�N�-��@�=���BJ1)@��1>�る1��R�%�K0�ax*ӂ5�|F���％���?[��&-����6mi%�[%�F��%�����(� �21":��Z���fb��O�A��]�[P����(݊�E�M]���b$g/EtB:�C��O���;������UKW������]�I\�>�=gqM�N���01��t���3�J�w���y�;�k��-�෢�����BFJ��#���D$'f#�:�x	��GȢLx�����Z�J�@W�������pCvdF��J���HF�ư�"�:����@痵�Y���I��w|�ag�X�'a�����ܳ�x���0���P�},��!*:�/�������z��i[s=y|[j��ѢF��j㏰�o��2l,���n�W�1�#�������֮�(�R~�G�����z���k�������v\����ǰ������=q<b�B�.O4?����������8w�?;�o��������8��y���a�m�'g�TX8�!,��J[wb�� a�t�)a#Q� +����Z���e�m�E[��)cܲ��=s3��Ω2�xf? ��U0/F暇��?�~�g�^c�}�z����=|Ͼ��mڌ���|�!�����kh'������nb������OP�j5��؉'�z�8��G{����Wp��_||�������,"��ߍpϽV�ok>�N�gKaak7+i��D�*�� <�x�,�CX2� $���Xz��g�ǢG��IX$o�)�=7~=f���q�p<!�uF��y��#3r��1�Ϗ�K�ңĜXb8A��]��'��b�[2\����񏫀91<;`91��q��H�LqJ�TBfA#��	�]�_WA�+�}�1�;K�ז�q�͎��[��Ű�.�}o�bdZ��尽eJ`[�b��V\�2z��T�Sz0#Jf��Y�SӐŘO�J���yD�\I0Q�����D.3���5<������-P���U}�E���2+,�H^�9��\Ix�q:���뙅.�yp>,�2��3� d��������{��eK
U7�Mg�.���N���K_�_������'?c'�?��=��jN��Yٸ��p݅�����^թ�p���D�W���-�z�1�;�æذi.^��s/���M"��:ɠZ��e�� �1��4����K���|.8��.İo~��a�MB���"Ҁ�`��L��,.#����q�7��D�*�X�{�T����W`21<5@�|��%j����9㘂{l0�2c,�p�E,�{�{����Ro9���q�e�����&w���f2c��1Ε#n�����,�$�bL򗡣�aB����io2e8i�xzd)���Ɵ	���<�Y��Yi@�2�{�\�:��.bX!�MF���[ZĆ��v�U,+f�z��E���~jh8f��ؐ_�pG�t��J�F��H*(E����S���6#4�A������\D&�".%!�aHJK�S�<���~�Ʀ��o�E���:�����L�J�p�\ｄ���o���gpE����ŝ�Z�+����͸z�Ο��o��ҒU�K��W�������,^�k�=��gY�B?���#p!#^$��Jz�����;A�,��)�0��0��x�Ѣ@l�a�7�>9�ᓽ��D�y'�j!I���;� T�ۅ7��o��>N�9�W��?�^���#oA�]�u�F��w��Uݣ��6���q���z:Z�t��Tښj��sO���b"��á}\�w�������!X�1vG���I5	iD�u��8�(*���je�yS����i�������Ul���Bo�..GR��d!3%rW o�f��-��[fY���7�YO�@d�6��:�u�30,Q�+�1��v|�4)�攰tH�Fv`��ĥc�x��`Ů����Z�:ڈ��^�������Y]W��Ë���^~�.�f���!�;��&'�~�]��/��F����?���������ȓsuCz�*}8�܆�_�P��4������]
�V
�<>2M��H�-��k
ªdxx5�_ð̗%d9�*M�=B�I�ٙ�\�W��g��aNoÿ�[-���C��gZ;��;�0љ v��L�֍vO��%x�d�/#O%��9���tC�v�7�9բC�9�LXJ���^mA�2�^����������4�z*3�W�Z���>��S��0��N��U�ZRC������4�L���dwI&&{db3Q�e�'_�6&J�]C&0�2T�q�ZҘ���g&��#&<N�qM�d7��Ga�g��8#1�>�>�z/��c����kB[���=�9.�z����Ĭ!��>'z?�ş���#���Rj�O��Q���
u\���'��g�'��/���ӟ��O��"��|O?�l��U��u�q�7�Ͼ��*�b�iNÇc�_��X�X�`�*"�qİ|G�E<7��H,��{�%�İS<o��0<%t%&�aXz���C���/%�WRL�+!LKN'��Hu���>����x-��!����/�|/�6%�	d;Bٞh���8W�^30���ɾ0Ez��_�)R�H�����n���a�cF�
�ឍ��wa�SC�[N�g61���#0�1:����t�/bX�G���cx4��a=��$�{:[�өS�n��a馇���a����Ű^����BX�BD�娆(a�I���oH�/�}�����Q֟�~\���˸�_�~"���<!v��g��v^5��6P���q��f^��q��'|���X�q=��JF@$���g8���[�ň{S;�KlE��LՊ][��;�Y5J�ڵ���A��Ai�XEk��s^<׹΋��}ߟ��<�yE��/�=�U����A[�������
�R͗w�q����Ӑp�ʻ�nƃI�lN�7�e���/�& p��{������q�T�1�XI�0�҅�f@��u���]���k�&jC-�ɭ�E��9Nkۇ�S��tVͧt}�j�!e�����<h%�g��Q���{%����^�<��[2L�FC9,�l����:ʤ���띝II1q�}��]l���������a�k�[���&�irG�H�oa`X��Hl�\�R``8^��.�@>����EK5���m�w?�)NZ�_�%~}r>5��rSLH�;���X[��i�'���(�]JN$�a�F$���9���PEoK�A�U/���]{�w����xؓI����C~'�����M������뾩���ל󽱏���>5l���'�7J)q��8~dB!����Aՠ���0��g�H
���c��	a��˘W�W�hr�b�kbKxm�i��ˆ=��=M���O8E�;]�,!�9�L�\@�����z���1��,n챉"=
L	����c@2��r�U�u�Bog�Ѣ �/#޻���|�;�c��Fә���s���4��g�WY�H��ף'fM\�i�y�?�H}"����Y�e�Y��=ֳ��cY}s)�#��#B��;}7�8�x/ �(���L%xP��0�@�'9�����:����y�|O7�OI8i��8Z��82��brc{�)6?�58T�Pr_c��I��;����_�>��i�	��T#m��X`K�6���[E�j\�X{�V�ǇC%fn#���B����Qe�?�,�������/Q�3A�����p��B��+��d��d���S��@��]���=��PG(��_�a��~i�ĭ�@qZ�-��_�DL�%hK�j�.H�=�4r������١��SQl�Z�Ρ[M#��@��;�����^���B��H����<�op���x�9q����� �5ߖ޴��0��ɺl|RIVn��u�N��C>�f�ܗ'��X��ORA�E�M��Ѕ��*_rq�.�g������LW�n�j���{��]���n,x��?���>YN��r�k ]�+���~}�s8�ބ���Ki����|�O-�zdi��^��k���V���I�<B�t�R������oO����2����%U���1���x��Է�`4���寝����#F1�v�<W֬ޒ� f:*�ٛz ru�]!N�BӲ��Q�>�Vx}2�m��"�v)d�,5)����|�T��q	Fwdv.���Xc��Ck�\��,���Y���׸Ad�|#��$-W�A�7��(H8[�=hVN>�����&�w�#á�A+�õ�������iW��W�>^�������b*���N"��`[�@ Y��Z�
�8����+Zdt���y�&�����a��?x�J8f|[�q���/ �N{25H��U�~P�	� 8<�v�L��]��V~�(`�ƑK2������=-.! ���q��</�L��՜��j�=�I����_`O�=�����㌸����i;-?��+(��%� ��l:)�LJ��W����՝zeG�l��g���}���u,[�J� ?j5�)���XW�?
�JZ����u.�A���v��b�җoK�l���#���	5ߕ"b�ql�/V�81	��?�EdN\}�y�R]��t��.3r'�/%u10�؅�y:���x����-5�n�|W3�;!�H'�����-!ذe.��	���H�50��ޯ�:(8�R ��I��~�y��)xF{d��˗\5����.�"
��#gGS�z��g}�{9�F)���_�+�6:�W�e ���h��6�RT�i�<�~��5���S�H�b��g��6��Ct�q��o�� �����6:Z����(�'ɧG>ҟ#�6Ze���]� $�Q� ���5@�.v �j����\��ʣ���,�׺�h^��Rd�;aO����|���`��{� �����7�pm*�?.��+x��}J��jЏ�䢒�p�*�v�hT��YN��{��e�X�\�?���K����Z`���c���U�S�Mߟ����8"<�1��i���F,�Vڐ'��J�|$�;����z)Z���A	���ܔ'�Aa�SWެ�b�~�k"p��-��JL\�/b3׾bvz���/$�s�i���#����nbW�Թ�H\<�����mS3Vv�`��?�I�x�o3奼���ˁ�:��B�/��QV<� W�jx�>pY5^��;�b�p�0��8e򭷞�����d���@�g��D2�<s?eCn<��Xx��&H]�^$�{pg�����䑤�A#6�do��E%~n%�D�+t'�k��Fl���#�S����8&=_L���=]%�n�*6�Q`Q��?�t��J�X��$�'�V|伛L?p��&���E�a&l�X�X"��B�޹t4"]Sr�d*+���漭7;��&���v������=��./�c�M;��Ү��Rf�Ѡ ��4��Y��ɰ�L��*�H,��y���ȼ5YtWW���#��<w�葞qZb�G���[i�j&'A,���By�L��� �F�������ׯ���1�1���g����Ļ�ڇ-{SU5a��%-��_�>T�߯\�<?�v\~�!
�j������3��j;�� ^����/���8��G�g���h\�FN��P�ϲ�G!\c����� �.�l�Y	FG�1'�w������<�I5C#��N���Ab|a<�����`Y�;)���s�<Y��5)g׋3�ɾ��h#����%ߣ/�eo�k����U�B*c�q�7F�>o�Ζ���(�7�F�%���P f����˃T(͒N�ĝ���C}j��~tΞ����U-pW�@�!s!����"'�9Hw)�.�W��ۡ8È�a�Id�t�i��%J��Qk���\�f��9��� S�z#ܚ��w5��t�A��Ny&�sFX���:It={�VU��`�k�����`u���\�գ'_����u���Ǒ#��#���:))�B>�MؒCa���"L�e�S��E��ѥ��ۈ���w֙�v'm���/~��E����� B�z����N�x~6�����6��ٵ�;��7���S2wA�%�^A�>A�������h$U�*61�{�xa�q������\"{��,R�(L����82NI�Y�?�(�F���b���|r�k��9��6s�/�8�+�^�4��ծ{��-��7�W��"i-��]���蔱N�b�h���H>E7+��39���I���|r-�"�1o��:��O�?_���h!P�F���������l��!Er�gW0��.�)�u	�T�N-���*>�rU�Ԅ�:��F��	6�D��3̹ٚ�^�8�H���װ����A�=\�d,�=�6	X��K%��>F����6c�����R����i�w��UL��V$��/qYrɣ��%U�P���Y���T����:)����#c�l��##Md��J�c��x�	b��
�r��S�=u(����.;O-�?���e������+�K�Y=���Iq�Z���#ߋ2bњh�<�]A�- F��=)�;M(%�NųfQy��!Ȅ��+p|�,E��aE�U:��&�6�d���:��|$l�����=�
?P��2JTQ8��_�pE��?;xCXN���z��"�Z���u�n#��a��iA�~N���3q�&�&t�q[��ͤ�LY}`��cM�Z0G��+�G#P����4��2SLN�ȣ����:��f��c�7+�l�@d��ΕK���ו渕E%m�u!��ǂ12��E<�z�J��uZ�F���w����4�c?���b��r?�Qq�u ?2�MϜo�Sw�f��JK6�~�L+�:�m8��Y�2��O��냿0��XϵN4��������N�U��^7ڕ�[Yy ���d��{}��?:�H|�-K?N���Q���)���W�JC�I�xlk�nn"t�*\�đ�I�{�.��Ĥ���Q�uP%��-�I��	HpL˻�_�-)Z������{�6��{lH�9wP����	���˝H3Ȓ2�k�%��\G�fP�;�U1�����O��/1���LuW���á�`3���U�g��&p�)������Q��rU���.j����?�s�?St����.!Q�k�;^��%�e�dpS��AҶ���1�(	�P�q�������*��4�7��,�À��IBJ_i��E��P���x���߃��l�g��h��'un��,�1�j��>��k��_?�	� ���=E8b�޷����8�Q>��ʁ��z
����tuԡ�Y/��&�@��ş�x3u�$G�_V��:�ͮ)���%�|����"mr���R�Ad�t`��Ҽ�i����I`� ����1=ZZ��r�H���#��>A�?������U}�8)�x&�=%*�������qu�з��b���8�� �\e�oi�M�+@�4>�2�.����kD��
d�2x�l(�^L��g3?b��K�kliy�4 ��<����t�Ek9=�O�V�^$lZ�}d�I}�i3�(_��G��d ����b��#�8<�GK��帣��F4O;y�Gu���wg�o��gZ�rah��FL�=�X�]7�X��ݥ��HyU��Qd��j|�խ����6�׊N<A�����+����ُV_�sڵ��wm�8p~)I�~v,%�V�"~g�1%IRv���'_�v���;+F?����q����|?��Q��ʕ���I�ʉ5���_����$F\4QR�<ze�h%�>S�-����f��[�mܘlz%&8�ƀ!Z��b�M1�������^��U-��n���1�ᤛ	?Z���s�B�0=m�2�KL�ۣ9�t(��[�F����CF��ګ^f�~�U�[�ޜ{̫������\k}/I���X���U�fK�A�:�]���"�:8j��&�$T�-��Ƞ+׃���*�u��m= U���*�|'���٩S��řT��!����Лe1�I��f�/a�L��G�>��z����Ւb����m�z�U�T�y]���ym�yv.i���F]K�T|]��1��Y|�������Y�SZ_��}f�g�'����(W�WԔmֲ���sTc�$���*�%y��$���,^ǯ��YC*�������l���4��pD�GEjWҖ~D>4-HOU}���l�#C����ϵW�}6�$�'t(��N�$��ɋ\����h5�e��:����e-BM!Z �؜q��ڔ�B���O��N�n&��#Qⷐ��Qm-�<j�Ԥ�~ng����Y
�`tq�˹BLwF�!�x��O�
A4CΞ�U��r35���*��<�C��zA���@Jے��6!�A-�ή�=ϯ�߽G>/\�[��j��\�y'����>�[�p�ԁ��F�OO*���>�I��� r�1]c
�u���u�V҂>o����/=��HX2��>��_.)�Ӽ�#���)��:� �WO(C��PO���ꍠI�R� ��ϼ��N�_�rg�<�j�F����:��Ʉ'l���BI� GD��P���!�@
k�x1�_*��"q�hzO!'7�A�6�9˳�3�eg4ͻ����O���A�:~���./���<G�⇷,{���M����rk�u9��Їz"	?���Dɗ�[��	N����g�V�-��!BO��'�.љ8���C�ϘM����Q�� _G cS�hL�C��s��_���M򻼏�V���jJ����c��懔Au�W�]�	��oH���h�Qb�y?g��QpW��c���
��L�hrR?�/�����
B��Gr��i"�Lb[Oq�Fv�n��bQ"PG�	i�Ҭ�L�@��7~�gE@�е���^��M�>8jY�"�&��������f����6l��*J��u;��Ǿ��T� J�6��|�nN��`B��{�u�a�,͐��&�����j,��]�����/Y�V�4���g\��.a#�OA�3�l~gi��Δ�G��ħ� �]�G���,-[C�dm8��R�a���m�~�/}�E�S�G6��x��[Fc
&�GvTۛ��~��=[3���yc3=,���I������(k����9���x1T� ���t��M�t}D��n�1�;촋�<��Rp^�ރ���^I��b�l [��<��>�!�����NZ�)�_=�/+�h}���֙���i2�-NqO�HD�Lƺ H�5��,�	�F�kk:��{gzԙ�?���E��ǞD��~�����g�%�������6�<wf]*��%�IQk�JZ�}�'C��2����0DZ���8��Ơ���*O#y��hF7�P�;l�MU���κ-���,�b��~�a)q=����SbV�>H�ӟT��_2�v��!��R�f�ِ��;T�چ|^5�H���_��m9~�H(�'�+N���щ�@�@}�������֣�*�,(����w��6܃��K��XJ��4h��݀Ki߬���a�2xb
(�1�6��W���*u�Fʫ@�P�*�S����e��Օ�X������d1�(�$�q�Be�o��ݳR��߽+�Ҽ}�a��f��9v�C�
gs��F�X���ЧS鮢�5�C�-��BO����V���̑��?ܻ"��2����?�ݹR̶x����뇩Z�H�j��ک�7 _$����V�?��D%��c���ա%#_���h��j|!�avĢ5�RD��A���X-���J%!^�]l��S�2�X:`��-nv��ɣ+����L�9�q��On&�g��6;C��f��u�6|�����N�n?^���-���
�+�:�D]W��K��2Ub������^�M��aV5$훧���A>��{x8&��2��j,��������pZ��~zͮ�臫7s�"�_�s-d��G��8�GG�:�[��J���Ω���5�c@>o���W#0�ߏ�#����)�ć$��>ǖ��X�0���f��f��_c{J>Gx�%h*&m�(�k,�QLƉq�4C��"~?HFĔ8��K��	��?�ғE�㒯�ɅM1)�`G�ۻ�۫�th���7`�C�Ӛ3���YЊ*F���+�:�:P�p.t4ٛ������o_��&Y�� j[bM�Y��С�$��{H0�Qwd�<r)�F��m���v!��y�XE��S5͵��4�阘��+1�YY�1i���ҿR�?��Z�Wn���e����T�5y�m� ��=��-���Y�`�(OZ�Z�	I�#���Ӯ҆Y�CU��hl>�W[^�g�?>���{�����aC�1FA�X����K/U;0�/�h0��JK��sM�g�!Op��0.�~ ��LRdQuN.���ڌN�t/G���\1(�W�@�-`WY�� '�4h�;Db�|�ty_v9�奋P~z��^I�O�>]6'Ԅl�إQ�K��ƃ�Is��w�L*�NH=(��<�>������,��Lmbk�T�,�q�w3�M=�(p!~$��r\��BX\i� ���z;��
��P<+M��=p�Bp�,�o���7wN��ǁ}�vFa�N_%�&��z#5��^Tu���e��9L #eGZ��0�`6��ez�����?���_�b��jT��*_�ڣ��2��$yW���v�X(�ky��!@N�M�(8�Yl��5����O�y+�H_���'\l}��D)fg�#�]$L�q�_��m��C��?#=z,��Ľ7��W�{elzg���Ƈ��{LD�%F�L����\����I���$oc8��vr�vY��lu��cix2[F�1��_���n9��+����+[��t��i�Ǜ4^=-��*�$��o9i��1dB;���K]���c�"�D��g�tvq�����b�m|�8����]7������������SFI���w�	IB����f�(ǣc�����՛�����Z�]��=D�*�۪y�CV��f0��j�9z�����-��;�2�� ��aa=�����h ���Iz�)�F pe^�
���e����� )��A<��.�G˄E�H}'�g��=a��WN_	R�иVUVsqlJ�?�qL�.�H@�}����͂�/�L�۬��y��f.o�.]�P}.K_r��h�aC>C�;Ay���nS㑴��w��d���8|:v��R,���={�� ѵ��+����Z~��q2s<� ��5Ώ��/������#�SJ�)��ݫ�`a+ rِe��o (��r��L����c��_��tU�k��E0����C��N'P���;�&Ɲ����'[�RJ������l��H!%�l|H��wR�XM>!���,n�BÅ-��&��ٯ��o��UC�S���?�(��	g^��~�<�a������(���U^�����4�R��h��Z���j��/NZ�)K*΀��N�b�{������/�I�P�_��KXƫ?���CZn�G���]���{5����掐^��!�'~�QzGƱ{�_vIV�#gw��9mr�}C��M���q��{I�Z
�)�f�d<Z���I~c+�V16�c��h��X���Fj��۟綢��+�C��3%�=5U���WM��F�͊v�����7(�=R-�b2ܩq`�$�̧�x"�q8�k���&͏��}��	{�J0�O^��[����wƦ�!!��}@�|V��!Y���0�>Lgw].E80���A=x��#Ov{d?�p������da�X��ˎ9ty }� �J}�Z^�1'Gu�( �3����7!�2�@5O�HA��!��Rh(P�k� ���&m�Ƽ]*bWG�࠘�6T�K�4���Pr8'�N�`p;l�R@KH�x��� �4~��h�@:�~q.`���gX7��?L�.���ly���H���)~b��'�z��T��w�/��lplX㺅~�����J:�~�p"��2BnuG��5.�Myж����%38��u���z#Y�p�����.�^'��D�nA �8 ������嚦-���b��CW�T��.�"���2q?�)��-�5"�G���Y x!�D5�!�M��T�A�W�s�`S�:R�#�o"]^6|��H�܏��!b��R"���b�aсB�Y�F�Obf�)�S��Z��o�<����m��dh#'�Wy�S~d�W	ȕ8�jV�w���m��~Й��J��t]���P�?�1T^*X��� �Q�ON�
Ү��k���V����9�A&���=9�ַ�;4�g�/I��D,�)�y��,����v�zh�����w�6O^$8���4�x�?��.~����'�b�d�kQ���[�8�.N�CR���!��~�f;q��6ղ+"�Y�8im�o�w���wC�X
�4_}E9,� �KĺIaW�.���u����n���2��^O�w����6}��t�!����F���E߈/�]�sJ�<0���$V�|���ĉ��P"^�iԚ�eG���{l�v:{n�S������GamF�y����>A�A2��q�.]Em ���E�HzH��"�%�iYwW�qz�f����6G��%����� �XR��-��+F[ݐx�b]�[������9D����G�,}�aT#3~F��	�B�*��6���,k�۽W���� ��B���w�J>�N>�Fg�S����%b���`$-��	����E�vz�/C���F�|�ӕE�'7O�vPĐ��¾l�oη�g@V�C�8q��'(��x|0.9�zP	��w�Cx�$��-��.k�Z�$����R��%; ����>qXO�0��ͱ�$��w��������͡�!�c�%��g�ցlL��u�x^{=%ăW�� Ǆc��e�� ��.����7ӮZB�}q*��D�F��;�kV<�F ��_%���
�sv^�N�� ��a�P�����W�ӍG�R�9�t����whM�PO�W�
`�c;��4y������&vqq��b�D�L2���F�e��Ğ|���Л.�e���z�Ϩ�W��w�(��?a��{�~8��f�t�����%;rό�O�!��&h 9��~��!��V��$v��x��R�T�_%A�ab 2V�x��U���%� �UOvE
>���==��C�f�䵷V�0Ҿ�rN��E�]!@��ay&�ecTQފ�_�"IUD۱h"���.E��[���/w�B�[��MҌ��M1���{�ӿ>�-�H2PZ�C�.-f^,R.Bf��Kz�$vn�੍��D�f(�xB>���̎�d������$��=M��t��q�d�:�b������	#�z�Homк�?	�7 4`ZY@�.h�Ƴ�0v�m#�z�Z�-zB�5A��S1����2,�8r�s�>'!���~4������|�jw!�%<�g���@�E�~�es�k���#���"u�P�=�˥g�ܪ�EvX_���s-���8���`<�	��`�G��SBii��@�VX���Y�����B'-��E?�[;q{��>:�F(l'���MAM�!��!(�Z�k������PwV��Y ��{h�Ds��=��{i�h�Ѩ�z
'��_Q�!���.�����L
&ǘ*�۾{D�k�6j�=r��b-Ċ#C���� e8C{�_^:�B'K���)��_k��D}6q�%t�c��Rc���TSr.CA��z��� e�ܚ�SB6�>ڎy ���C�\e/f�2jI̝�kۼJ�� "h�������J/����n��I���(I�F�Y���=�i�]x�Nc��%d�(�!%w����<	J�����/��Ѱ:4c�����A�N0r����K|�2��T���Sd+�S�	���6m� }���[H�D��o����!!/V����G��l͟�p���-���q_A���,�|��)ح�Hʿ�~�� @�ϧ	սl���ѿ���.��]���nO����A
�.���,���׼�I8�f2��-VR�L�������-KK���q=92{�N� �g��)��w���E<[�e>i�w�ٽC��RVĕ���)]A��ו���J�u2���ވ[8�,}���p��\���������Њ��:iey~'��y�찕��/��y���X2}�z�4��/�S�����W�x�b{KϠ5��J�3�Jdu�s9U�#*��2�A$=To�H���`��Y?!��V�ߩ�����j�������?қ�N?�<�+�M�[���1]v%�UD�����n��G|q$��?5�����w��.��^�/�c�]إC}̘�MZ�J'��&6(H(��G���?]
��7f]��S�O�X��7��#����<tg�;�&��Q"�;'��ǻM~�FO@y����_��
H+��oZ���@y�=to��Z� ��&p�6~G�����d

rz�w.0�#� �c����Zȓ��-7W`��P�`�}�+?[�Гfϰ��hA����1�..��%��A�Q׷��7�/�� Ӹfn�_��-$�����/���ۊb��:0G�2��@q٩�4U`E�!��p��RE��t�#�}�5��. ����\��� �(
���~�YI�,�1` ����*6P�t�\M.��^
&�������S�b���*�+@��1J�X݄t��{"���4"��Z�^7�P�n-�h��rZ�U�/����O�؋W�9pj���wV���Z��,G2�T��M�x�}��yČb����/Ka�=\0r�sņ�|�El՟�׍���F�~'ő��6�	���nB� S �!IV�pw2nZ=�ۭ:qb��WN�w�vj��E�D�T�&J�X�q75�֔��̗�2VQЛ�n0���6�i�w6q�*=�UЩ��z��Ll������ހ��2`	6�wPC�G,�-�\:�♫�T��d!+A�B��1�#���WR�r��\�eX��Xb��W�6��LJ����])��s܌�O;�B�'e�Hre��;�u`&�"e�?^f���D�R��j�%�5_!j ��4/�3#p��I�/ �����&�u`(��R��e�du,�1\\�Ju &L 2��Siq���Ev-��v}�r��k��v.���!�~�Ό]��/�K����E�~��b�<<R�ֿ�HWx��UwK��<�?Z/� !�[%dx4;�=em���b![���\�������|>������{�d4��ގ<��a�]!����3��9�ٜ仢�B%��̢�<#%B�v�>mn��f�[�A�M��#9FO�!� 1���{�p�؃>F�������"���(�e|��^�_��?����Þ9��_��&�o�<+�ʵ�C�z>Q����/V4 d�A`�W(����k�1-�e����%I([�?�Ԙ�u����1^5m��ܑ���`�Ki���{G�u���\����2m8A�_EO�v/�`�6��ן]��G5���d[�LҸaE���#}�o�s���絟0a����Bނ�S?��=;�� �x���j�O��ţ�B��E�u�/�kO��(� K�a�u�s$�?$�����-q�H~l��T�JЂ�}\6bԢ��P��(�V~&ܝ2����,�x��TƤ�!��8�!���G#������πL�j�D�ܣ��H7ݖ!��i�7�q"���l�4?�.=�Qv�4y�h���Nr䫳C9Nh*}��m�;f�}��ƕD�$�̹�l5�oM�O���o�^�"5;@.��r��0�֌�,P�ƞ	 ��Ŷ|q���$Z^Y%朚q�X�8�+O�֨q��F��җ�ZC�?x٧6-ͮ��bdLT��J��L�Jt�N���#J��XJ�]Y좎4��K܎f�L֛�K���}}9V�C��/]������_]�ϟ'--�M�jȦ p���0���3�������k}�A�Y�jD?�nE�-��co��	)�pq�h�Ol�H>K�	a��T����;N�X'㕜r�ƌ1}�a|�\N��J
�.?�9Z�Z�Y�4ئXr�������ς�H���-��9:�c����k���+��H;����^���g�9%d|2����A��:�'�1h��Nf�e[RH�CY���*�}���6é�R��k�wl��V�s�_E�R=ݛW�͔��x�<9f���]A���k�\I��}kZ|<��i�;�aŨ�����x.,A+F�+��=��v�a������/� ��
���1T�-n���&�rZr)Q:<˵/��Òc�M���:����͆�i��(��\J�u�u�9��0��ݞ
W�{�� ���l˒�?p�3��:����}��MP�.����=�D�G�k�ڧto����y ��b/�q^�Q1��xE�F_�ŔŊ�M��$��IR��L68�1�:��}F��8i"��.�D���u�Q1��c�z࿣�fl�/���f?��M�՝��o!b�0b�|]&p�և�>��Vn�t�Qv���_���_��H%�X>�d�^����*��u��n1-�GHZ��:.n�l��S�J�*�f�M,j㚓اX2��N�[�����>Eu�t���%�gƋ�w�G .�6�G'�/�J.�o@WIl����jRxm�c��A����y���'\}�}����P~�F���}�u���u�CMA��9��������m���Z81JP��ܦ�aX�0Z���FSǸ��"��)�N�����O��F�_��sl3�d�8�#g�
S�"?#�l��XA��\=_z�F�\;:�nQ�-")q��d���`���-�sy��6`�ày,��!q2���]	�LH��4e{��$��$0��x��{xi�ֵ���Syr�K+��+/H!�1��h�}Ӡ��W����y`p���OߕiY�%��$
[�����lб@1.u�eN�:��f#̊�����lR�N�/o<-�K�K���bV=�V����%�E�z��!aāI�p�䤾f���߲5F����p���&;i��h�h_֋�P�z���t�_P���gpE{8B��	ۻ��c���E��lO�*�1@}�C���?���Ƀ�`"2�@Bo����ِ����`:- �w��$�I�����G<(*5�H����VѰ�Ǹ���;��i@���(�@:LIއ��B�Z*ߓ��(��̴
�f֖O�^��_�x=4}�:����6=��[o#Q��U�]�HLA;�y�d��Q�7�������	9�R���'\'q,�vh(/�Uض��YN��]��m���Ǘ���"�)��S+���-0��]�d��y����/mG���W�͆��V�/:��t�=�ĵ�:.LjQο�]��I�ۃ�?�����dCs�;DH�҈�e�i��$�ޙ��2��
'$=ĠO��>1�O���/[hO�"�@.ƻn�?{�ῼV�GVJ����q�?�l~O1jk���{��.��������u;�n&��]��f�$i %& Ց��)��B���Ґ�Zr�#�q���� �8+`���@��k+:I\�:(A|D�(�Q�����������~L���@x��Q�5ˌ Ԙ�����3�ƈH���RH�R�јľ�f�A��󟆈a�#Q��i�F�3�a5���_�s�x-u%���` ~u@�Y�/,t���M����]p��2%~<�����}D�Xb"���V�I~��3߂�O���Hv[A(m�޴l<���U2c�[�m��m���=�2O֘�[:D��)�����K)b�c��w��|q�	�R:6[�X7I�Ez�ZF����<�с9���ޑ`Eӎ%<�3���](Z��aj���~h��ֆ\{QG�ʫ��F�Z{~qJ��#�f!L����A�7VfbZ��7�y�uGvԔ+�`:�Ҥ�e���R�.S���}�8�ap�O��E$&s��<堻�X��KGI��J�`�3PҮ`�?`�N�`���� �^�1���ED�*�-u�J	gٶ�2�q?dhSG��d9	�]�.��\��O�ǗKٝ�Z������f�cO����(��"C��Q7.�)��J�������<8d��������AޔO��hP�̓k����*���a�mV�ߗMϨ�\[2e{n�O~��Yj�̕���D���jN$J����p���ͮV�
���ɷ�� ��3ey����:��ʥ 08ʬ΃/`��^ӻ���� x# ŋ�9�u}��U����(�knC?v�`�-�KD�|$6K��ĊA$��7�S�Lϗ����%��ZO��<Q�ug��+�>앖[��&-͖1Z󫄪�ߙ�Ԛ���mG�m�>je�+����;��H�xrG����Jؼ�C.=6�Wi��˶��|�6���š�_-��?dH:v��*@�!��ݑC{�9˳���� �%���PR -|^x��m����#�@B�Ԡߌ��IO�?����'���l+q�z�rPn�u�`|�+ڠ]P�4�	n���u��΁�1�jTH�L��k؛�N�xHB`<�=̩��+b�r��?^Ú�5�4L����<��g��k]���k��+��X�{�!4��g�y�v�m�x�-C�yCctThci&����>��ѻZ��~I�����3�఻ʜ��يkm��J��͛P��i#� �����zP�F�7Nˆ���[��Ô���'QMOw��-�8�\�uL�y��"yO8C���]�L�˖��y��d�`+���x��x�>�Ǹ�����'1�ԩan�j���������w�?;��.q!(��"���Q�\�*���NR��Z�������R�����N���|���J[KOb�]$gf�ei�m���w��}�{�f��$��[�.b�zq\�'�r��OAt��ޔZ�q�U(����
�WS�I���8������9�����˷���'�"��5Cel0�^���t��@�B��5s١Jb�9�ЍV��OB��M��ͧG7G��IܙeC���N����躣���?!F�WbW��l�V�ԎQZ+>��;�,j�j��hkoT)�Vk��+6��|�ܿ��s���>����9O�o`�㎕' a�pk;!�e=t�uħ���/F}�M��>�RА�@�ۚ����|A�N!|ЎŌ"'K�F�:"�k�k"x�(�2{Q�%�%�<,�N���y���(��Z�'�2�D��xt5H�o�?�E�yV�e)���V��0r2�'�i��cH��ԓ��������Ə�E��M�f7+,wb(:>{�{^bS�����k#}��j��m�?�/�bš��3�0��$�U�d���~�b�n�;K%�aa�`����\M��Ʋ��w^�)/՟og�7ձXgvj����:Ypu�(4ks,��[*x`p��w6[������u�Զb|��8�{�KK�߆��7z�֕�|l�¸V)�]���EeCYq}��	~�++y'±lByc֎d��fcW.Uuq���F�DN��<}�\9\�����4�P7|0��8~�o��nw���V��n�H�	H���i6����P�An�� ���d�ZU��'X6���MВ۟��/qRѽ.��phiy�v)��	��\�n��O�o�\�_��/о���?Kc%ހ =�w,��s`U�d���r�lS���;�ۻ�P�a�m�Dя�'��C�xb Fd��n�'�'nT.��A��-A|����G��v(��z�E�(g@�I'��<@�Gl���������L��Y�\���#�}5�����Es.ꗡt����]��x��T?��ӬgHYS��j����SL��!t1{Y{5l��1��c���`�'� )L��趃Y<?4S�}1��f�Ւ�Qg�X��֊����gK���k����2PGa �Hָ_|��^N�z"����fu���s��ՆW����������1��~���[��*�QS�c��Ҝ$�bd�N՗ 9o�k����g}�gAL���t�m�V���޻/*����;�yp�v�p��Q�>�����d"q��H��inS�����L\���L� ��X4Ȼ�U޼��qbV-�O{����o�=�j� �c%8�;-|�~��$�hr'��u���͋�e���㢵M�]��yv`H&ģ�t��eccŹ)|9�-�L���$w�����N�49
u���l��R���7��I�^��χ����� x�����o��~�p���\3�UFE�R���)������xsh�W'�;���0��a��Z���bc���T�����-+�rZ�'8��m���%^��*���c��d�d�?��*���:�G�'�&w�?��*���I��T��L���|�3�8���ft�ȈʘO���i���@�*G|�}r/��O4�&h�j�X�Z����%�mqh��u5���Lj�l�hC������s�Q�&D�wg9g�562�|�DA~�o7X-y{*�E���C�#��sB��h=���~�i�ňg7P.����el��e�D�@��Yh��h�R���eF�Rt��9�~�x�S���/E�F��4��P=i����Ќ�җ;ZmW�M�s4;���љ�4�p�?��&>�G0�c�͚� ���J�[,�y+p��T>�b ��/	EI
�1?b"/�vK@��GX>��X�)"��#,��A�v����1����ٚ���=N�P���)�53�՚=��fk{��.k�`U!��l��iP� ;u�׃\�_4nRi�#��4����P�6�v2�r9�K�(���mw���
��$#u3҉܄kp-4\���F���x��U���V��=��H�e ���Ч���gIM�I�b�7b�/�6�����y�P#�ͣ�E����tT�3��i'���'��
X��s���ic��t�D���v�'��KBnM���]��_��k��QȵmN��B����	�_M��k���tqs�<�J�.@ǲ���WY5�����E�fۙ�:U��[�DF���?��\�wZ^|l����\�ԥ����|4���w�11'��]�G�MY[�t�e�Kq:v��i��ƅ�LVh�^�	�u]�-tC5׽5b���<�ԁ���U"s�����eO����yG	-�n�
���x�Z�����۱;\>���a���I0� h�p�v�S���N>k�h��v�$�5ތ+bm��V���&�|���R�d���+��ޣ��i2�S�$�|���jW\�vF�����l?�+��*�-B{��XA9�ȑ�10M����<pn��E�r��G��ʇc��(�~�%S��u ��y,ӭ�c�G%ڡ�Zzv�@�Xr\#��ǐ�vhv�e�e��5���"OD�zu�3��"L%���ֲ� l֕�|r"��h�� Nj�x��"�c���|+�|Q��+f�O��J)gu/����?8=9�4p�ej9���
8��sE�dsC3�g�N6��.���d�J�������Bv�'�'�������'#�C@����P��ڰ���a�hBw�6������_�Qp�Z��$��,r ��|���>̠�{Q���k*����'�����ɠ�c�Uj�3����PR�-�_'�Pfv���S�4���L���,$�eV������@=<o>�;$A[/��ߥC=^��{���ފ�����k�Ũ0}�i�tUS�qɀ8� ��=&�����pŢ\�ߔ;�-�Z��9�$o�+H�ѾdO��qifF=k�r�da; O晿4ꩅG��#������3�|a1�!6�P-�@�8�5bE��X�����8�s��Fd�#�Y����n;�	���	��0�v�P_��!��J�V���=<(���-���c�U(�5���/�x`���\w|�'� (�R�������=b���k�Q/\��b�|-{8�:�`Ih� �ϺsE~_�}G�K��d�$7����ff)���J@�_�|�
�돕��DD��;'�խ�=�_�������B@=k�ހ�V��LcOt��)�!"�Z��oB;���Z%��P�{��l=��m ��m������6�����N}�L%����&f�]:�i�����O-ӹ6���ʮ�o�mm?�[��B��ehS�Mc����]��g�S��^�V4�S������E����z�M����o�C��kצ�����_�τ����s���+0�k,B�8��%&p�=X�a�_X�Q�c
6e�����j�h5�`Va���O�����e
妑�`2ک�~:�?#ӯ���3B`��]�����K�[����B�[�O�r|9J���/��R�E�ͥ�1N	�����!{����c�C���b�5�~�����fR�Nz�2��(�"i:�����ʠ�S���ݝ�X��������"ZT�)^��Zr�	NtQ�zu�&~���?����VAE��cc�� uE?;ޘ�w��+ZM;��7	��^�kx�����a,.�<��\�$��$�7,P� �c	1ܿ�Z�*(<iX:Mqǚ���T#��MG���(bo�I9jj�3�O#&�C>�B�����\��ܹ��`�[h���|��s��BX�~I��	����7L�s�!�������LdQN��Ќ
��$������H����'`�eƒT)���[h/f9��v5��Nd����6y īr#�o� 6�4ͬ8e�'4�<�J��ўq���g�Η��`}�&�y+7�*�����Ӈ��I�����(�<�ȎC�r��b�^�sl,f5r�.~��S�x��vЙ�����В<Pq�n͠@�aLc�HZ�k�	1�u�d$�C�7�t�1jɝ�\�Ee:�m�ڡ����!9q��d�ۼn]D>���0d�94�I>�Ȋ��d��F��"�-���i��`�	H��7���E��2 �yleH��?첵�ȯ3���8��ږ/���,_���s��o�3�����v��.��é�IըW�1��T�m0���}��8��zP��a|T(���~����l	HtЯ�'�k��M����5S�O���<S�9�F��h���6��9�S��=B/.�D �&�S��#��֥�Q�7�sIɝ��xAe��I5;�T��}�I����d�P ��+a��9�����~�Mg�UE���t���֟-�l߽T���JW�v,�;U�K�<q�/1`
�Md��?:�{����>]��0{Sp�cb�{��a�t����R	�O7� `iؐ<�ku��Ͻ\�/�+樎b�ā�+�;��6��W1sb�
����E1.�5H��D�D���@J��V�B��O[h����o����W_C%�*��9�5����כ�S����@@�￣��ӆSb �"��ZL�%�o�Ut�����?ɵ:�	ot��u�������_��ay-Q ��pʈ�~	)�wa��<8J<hͳ%�tN�_3�BB��&����V��>�lP����όe}�q��ب��������1���?������}s��}B�"���äR�]5�b�9��Ҙ!�9J�a�p�Z�<��4������z���ү����W5SO����qj�8�U�I���ǾWw��E�=,(:�q�K��Q��{�5.2MS�'�/�p� ^�3m��-���k[�|��g�g���kNL�p�hfq�>�H�͍0d�P�o��V�
(�ZH4�Q��$>��*�(���n1Vv�l�7v�z7�wD�$ql��TAN���P���pN Y<��=�����g$a����n����sg�*`tę��y��,���Qa� ��c��}V�`�<�o�f����%U=ܾ)�� ҳ�����2g�qd�#�A[��Z�2G%�c�\] {a�n�!����	�N�������%NNV��wm]����d�0Ǜ���Q���&2۸s�r.B'j��V]x��9��I�Avt�+~OI��­�~g�_�� r��h�=�;5�v�{.�E�+w;N���7��5��*3�x�����s�Z�(&L�O6��C�sMϲ����v>����MdV�S��/掬���w�+eE���ye�{�)�'��T�"#3�z5�0���(��G��&�D�A$�[��Ź�h/��Vł��):k�G
� Lq�ܐ$jxNT��Gf�� �l���z�ȓ�mk���-���m�gԯ;Ь�c��3�b�o|�.V����e��3���SĿ:<�v�/��n��g��§$��,>���6��|��tIŨ̒k��878��
�bٻ?�z��m�%�0h����ĕ��J����/��0�!�pp/92�$3g�k�B�-gu9~��֔�_�>�Bc~�vO����nD��i͂�;�U�� �G��T�h��)_H-����J42��\?!�\�B�����"���S���:�
�
]��V�
! j���T���ߵ.�����R�A�%�ϲ��}.ʑ�^�/2tj#��^qM�}2��ך���%���m��3�%��T�7=�ޗ�E#�Xc51�B�k������� �X^���}��	����A:��e�k��b�{|�s7�>F�e�06��_y&al�["Ml�Vp�dx,tC��"�D�ߗ@��(��}V!�v����i�ٻ�5�-	pr�s�=ͼȈ�z�Udҽ�!���=9[������"zL�g*f�������Sf�@cχ�Qdʣ~�I�R������{{5��7��V�����R�0Ư��K��
`f��vR��si�(���/��;5���Y]RI� ﭼO�Z)�A�۲���M�jRn�_z!b�,�O̴�^�O���s*�0�z_���!���jr^߀	Y�׳�1O����t�*�A�i�"��)�/B�f�(�1>�@�N�\"��c}�[e���b~���������d��P�����G;D�=	)��ISق�,��r�p��#$Y�!�\р�_YE��1}���Ѡz&R����� �S]�Ay���sI�
яGtU��G7�io�����+����KSJT��+q$�sЂA�=$;#�F��v��Iq�]�#�mލ�.��Qҳa�g}��-�k��P2w��o�i�ɷR�h(��ɺ������*��Cm����"lT����Y��z��^���5����{e����p`�e�$a��K�z^d��'c�VB�ǔ�� Uɗ�XP���h����,Fc!$1��LV6����Y���I�1K1�Y�u�3oӌ�SNʚ�	�R�q�P�`5$w�)��Ǽ��3Ѷ�������9�U����ň-����c�`�9qu!��@Y��+�:�V�D�n�*�R\j��"��d��W�Vn�ځ#L;���"���T�NX�8�)k�8���}�m��jpg�zˉl~��YoI��i8�k��0��L����̓���نEJΪo��[�������(Ǩ��.i	R^�3M� �wS�3�D�"���c�����;����+g�uva�y�u�������ˣ��ˋcv������(� �'�T�*k����f�ڗ���ٚ�|�S��x�~p~#SF���� �7F獆���N<mkV�t�V]_���������0Ϊ���^P���z���-o��?[W��.Jy��%���M������h�1�}->�d���K����th��R�s�������orG�6c�&�2�=|�����h��F���]�jV��]�I��vA������?b���%�8�`^��*�w�	��av�3��.���0��'a*G��y���t_v�dQH.^Ha�Ǎ��\Y����8��4����7��2���2��>g=3lz���������5���m�3�HƊE��.�`-h��ge&�SI[w�����o�J]\���݋﫦����|N�h�+5�m�i9wڄ�$�˽�;x���gٙ�PČ�=�|2�>���B:�YN�� �.��,��;����7c�¿rޫ�&����:��p�^�A�������� rSBm�u�'��U��7�>��F&/���bK�C��G��Y$��ZL��Y�x3_%B;~ʤB��0�>c�o�dU��1�w7D�5^~I�ɂ�KOg���)���wǳv?����'�{�5H�֔��.ʚO�
�L��&N���=�������k?~��fR"-�Jt��"�
�'�}%�M�We�]E2>������ ���r�E'��>h |$�@�<���XW��&��3�&Y~f������I�P^iY���k�En�����]}7�Q���5z��}��%����G��o�-��0~��������C5�������3y��@ΝZ 0g�+���-ٿw^T=<=���t��{n�-���+� ���Ѓ��"���Q����
��d�n�����8��)>�٩�ڰ���$TI�Ll�������89���������M;׋r����P������'��Oh���p>�"���*N\�2MR69K�\�Uc
ح����h�u�I�����t��������W}�:%����L+D��ŭX*��Fx�~)  k��Sp����frL�b���)�_�o�)lX���{Z�����C��5�Cώ��b�h_��}@����A]�b����pf�2,��<�n�kk/��q���%�:$�{�.��[[J�ݝ����&
&���W��/��%6����?]`��ڝ���<��Km�Ɍ:���/�t���=�@i�eT�&WA���F�^���#���av�E��� ��gX���h����#�[..݁�{:Å��D����)í�������Z��ɸ�z�9¯�X�N�N��7�	���Z����v�����w*�Z/�N 8zl�bW|��Q�^v�$=ԕ5i��=�h����0��ȁ�+��' ���j�g����!E�At�TԨ����kQ�B��zyW�׉�?��l��{�Ht��-���Yo��Bs{�?b9xNZїJσ�p�?������r��>{|7�#��̭+�1<'�FB:LL��6ұ�:��hl�~��k����2<�p�j�>���Ʉ�o|�1cTq#�,��k�IZ��>h���S�Ԓu|��S�����FF�N�/(��%Z�N���H��bO`z������M��C��_uT+��}/�i���<��[ȢWn�G\cLhWD��ɯ}�1��k�uS�a}��U���� �KP�0:S������V{"�?Vo�Lc�Z�cZ�*�={5޶�����a�r���Kٽ���~���>��R����[���_jh�~&+�z߂㰊���4���}<�J ܲ��D.Y�]a����YA-�zǌb��_r��� �c��+�zp���=P��c ��A`{�T�J٠p�EG�C���$J��钵�A��x�j�O-���:/.��zӅ���=��*�}.�u�f���lKj\�\�U���Y�%F�F����
o�>kw��觬Ƣ"�s�P-�Y=K\�
#�M��(�Y�Â����`��r2�J�	�C�+�Öu�ZJ��Y7�тO���)k��5���|� $.��J�ts�k��컉�Mkn�I��A��`һ�W�vt6��m��S�/��k���â೙���RY��j��0WJ�|zN����+��W����S��|ȕ%L��Ƿ�Sv_���.��-�_$P��e��㾎�����7��ܯ�`A��
���o�VT�[l*U�(瘔�s�6n������5���qeH]AG��T1�`�S��%�J��}���3���{np�L7����%"�=��X$#=���+�v@�6���lUȂL��ttlxs\�gUs�YBp��=���NՑ�^[�O�A� ?z\0%�@A�Z����a��N����E@��6�:�~jն��ÆV�>��kO�0�m�"	��Kf)x��	ڸi	�N%��{�\�F2suҘ6�����+z!�y7�B����̃|7�/d��X�T?���A����p��G���`gx��+�����/�ݐ��A�YX@{y1ٜ�����\�����gC�+���A�G*-囻��N'J1_��k)E��������y�mؤ�����P�vu��G�n��U+�%�3�'V-�/v1Q΁;�����b��9��?�!2�����,���uO�&��ba����"�_PQr��冲|��M�kk�Jڻ�g^O8Y~3�B[����&ۅ��[�X�@�QqW�!r�-�n�خ�M4)N�V^��9�c��k�T��\��F�'��\����8\�鲔�"�������L����(&TBZ
#���ǪЀ���ws+���)��'cK����M����/%�%?�R.��c�>q��%Mzgo�������!��A�=d���ۮ��O3+>��8�52�����\w�W��Y�H���?b�w�نu=!��;Mm,���wQ���	��*�S\�'B��l=0��w�'
�Y*�bTq,�"���yЈ &o9v�꯵3Dϛl��J(q=�O%=4�
G�D���7~m6�[>�+!�QJ#����˧eHt����y���|9�gH�5Q�,�1���v��h@&O��-��t�Kp���1���ے��������$���a��!�y��΂��M��Rb�)�jmw�� SA9�����B\�㽻��s�Eǹ�b�Ҿ)��Ub�z�+q�}�+ϥ��lN��^�y���4�G������}b*#Q�O�N[���CsP��qA2ү�+��qaH�� 9��j���	�=8�J�Bʓ	�}��m��i���9,�t� �ٹ����-0�yؗcN%ӟ��<%�r&��Eck�剰b����Z+��g$-�� ���pÐk�����/
�Vbc(~F�����Kh�hJ�H�:���i`]�����օ��W����Ō�MvjL��< H�뚰�U�1Uf��R�z�i{@�³w������z���ˋ����5�˚[�НC%��|:G%?3��b��s�d�����d��+Y�C�'D�+�c�'�q�A:&�Ϡ*8��.S
Z-�1�u��T��bO����
�`�g9�@]�p'MR�6r;�P_��y	�xU���v���}�1���k�	�7S�'��b�ڴ�-˂�D��xh��?w�������'�c^���e�S薸�!��\��jBA-(d4:v����o�Kj��ߋ�A�[����i"+*oY��R����t���$�	����������z���M�p��C�Yt�����KP0��^F�W�!��{�s������&�0�4�&Ϩ�-�kK��m�d�Cr�.W{�
����fK�C�ye*�a�p���ǾنKe1�g`��<��v�.�Bp~��T�� ��C��F�G�Kz]�o�5�XC�H{�qy��Z,=������Q�+,m�"*`3lܥ�T9"$�k�Ќ1�=۞����&Պj"�SZ�/�z��[����oI>�u{���/Y�"X1����Q����*i�a��۲iz�Wn�
�u��a�i�c��k�\��g���ft>~�/'�i�;U�}�D�R����r��#��&1i�T���͇z(����b`�5C�U��0F:8q�{�0E����Y��=�;�'��D� s��d2�3Iw'�-���u�
P��A�ݔ�َ$�`Ĥ�uZ�Ձ���a��F.���ҙDY����~��SJ��#�_`�Yk�9({%�aJ��$>�?�r����
T���x� �������;)YQ���!J;��fɔ�%?��|Ȟ����'�� ��E�bb2A��Z��،I!��h�?f�4|�cІz�@��<�qz&y���z��G���7��cb�T|�d�l��e�Y,S����KB4�!���B�
#'nl���w[ң�y�ɠ���p�3]�mհ��&5B�&f��C&�������4=�=��e��`�F<Y��#槂18U�6e��� .l�a�> )�����ӝ�#H��uG�^�}�Y@b�H�(?L�����9ѣj���j�ȧ(����/����i��R�l������Hlp�v��ta�P�&�f��^�Y���##Dc	�f��xD��1�y���R�f��n�@���$�B`�f5���8-I���� ��o[2��3].�X�I�~��$�,C�/����N����G鵏�J�\��n��v�|��L�L	�0+jxQK�:�Lƒ㟿ɋ��%t��O NU<�̮tt!��ZӁA��Y<;���l��+{Yk��'�ZB�`��ρ��ŕ�ͶTe��f���a���}/NC����
j��+��樂a�ŋ����l{!^�zS*a]Q��>HD���qGs��k[N����y��ꨴF��8fcK���]l7U-<:�S��6pt�n��/�����!/ǚ�U�uvDn��Z���Hǩe����1�W�x��~�(#GZ�L��p�~���"��5����[��vw�jK/2I�A��g�iԹ�>4��@RB�. n3F��~�ײ ʓ��U���!Oa	�����v�
����a��v�T�&��/ԊvJ����^N�@9J���,C�r3o���X)�Q�=�p��ɯ:�B7�?�/����e��y8u,1��Rta���#�
.VJ�D
��#���� �� YJ��O$I�ZDC��#���7cU��G|ԥ4�BɌOM�~��触z>������ХQ.�6��u�.=�`����G�:�S~���z(��C���5'x���1��X��{�s�k���ߟ�x*���H�O����(JS>���\���*tW�����+��(�y��x�$lֺq��-��?vv\Ll_����	� �j��ۿDE��@_	c��8=��!֠�Da��nN\���O�$�_w��"!��pp�,���&�>4_�̋�vd+������92{�*������Z7Ƌ
W	�Bq����"��Ă�C�hau ��9�5� C}�����J���ل�jvK�r[�ִ����x*| ř�a����	p�
�}l�Gr͆�	e�0Q����ᳮ]D
Sg4e!�$O�]=�-�s^h���%e5�:|Zޔ���mC02C�P(�(u��D���}}�Q<��q��4�-��۞�h��_U�IX���)g���P.��{5�����&X�x	-�	��O�Nm�țKts0?R/&:�c3��)���ɒ�Թ���WxyE���j=�������m�!!�O�4'�s���e�cj��+�`Q��B�Aa7֞5	�g����z~uOrٺ�X���I}2�<��`�*���`Р�H<��4��֚�5_E����̔�����`��s<��n:[�)��_�M�K:�h�ہ�v>t�[9����J��&��襓X+��1n(2�V��l���sd��>��tUX�-�l� �M��XR�%^��/�˄yJ5�^^��+��S��1����_�<�KGx������If�$`V7�o��U���s�QRa:ȯ�t�[ضO��D�S�����%+���Ί�����hN�z�FI/L���}�*>�3�)/R9��4��b��,Jm�#��2�B���З���ғ�и�M�~K�Nw�S
�R�ӋGzb����؇ZW�NJG�HA���t��/��%�����]�Ҍ�⩰���mc�Gfz}�f4n�d�w;�W���%������iG�a��qstm׿x�Q��ހ��~���9?�����Sq�9˥�Բ�����_��׼�+�c}�to��H�p��=�
���**��A�N���3��j��j� d�wI\��E�=J'�XA����$v��훟�`�>U��9�{�?�s�Տj�$�?神x��ӜD�"�>lN�rM��jL���6� �8e�eL�����_�|e7m-S"ls����O�9��W��8�ܨ����_-���{�>,A��C�r(��]�3#k�>ҘnF�&=#��A�꫁���Ⱦig�\k�Ɯ꿭\�̱�e�'@�	���?��q�ٽA*G���0�h�j���&p6c��oq��B�ؼ���w�ggb�]�e�� f$�(�f�SZVth9�C�@"��E޹��y�x1�r=D��޴!�����[����v:]�gj��N�]Z۹Ԋ'�耐��U��Y���m�X��:܍F[p �ԓ��أ��m�P��fG�o؆�^�lM3T�HM�����abPYETF�8f�*__`w5�W���)0��-q�������f*Cq�C��xT�8�PT�4���� W�G]�C��X�|A��
�>[~��l?����T��.D|燵e ��A���U��s� {��p��̯�ߘ���<�Ÿ����8	��n y`ϥY��l?����$�$���8�2|+�-���z�%3m5���a�ʎ�b�5N�?���.�n~��O�5L�F��W�	�K{߆U��5_^�7&",S���\��N��hf�2RfزG'�%�̜�t�lY.��l�k+_������;��Q��񾑲�գ�H|�rq�Fz���]����!(󣮃m@�u��T:e�4kbP���I���4�����+;JY&�wOJ=(�T�މ�I������X��MB<!�my����K�+e��)p3eA���/�6i��*��6r��p��6����jz��A��m�	���J2��v±]��0���Z=�r,����Xb�q-�k[\T/��j��鄱aۆN/PvH&��n�}[�kB�#iY{H�n��7�ϳ�ZN����u~�Ҍ7���d�g�J�d��	��&�c��G�$z���m�_כY�k�tV�Ts]�����j"�\ �N���g)�Ձ����g跧��z��޹}���h�rUt���j��K�^�Q�?���:�k���^��,zM�A������Aq��y�x4��9��x~�"$|�lKw����!�\������Y�m����y�n��A���"古s����7���>kJ6�C��Z��X��8��P��CV��f��-��?�M�~�����`S��W D-*u=��{Ɗi���� �6�&��!�sC�g���Q,�)�>-�6�:��6|���RQ���b)��T�c�����;)+<�!B���Te��^!m��Y���9��6�Y�'������hP����n�śhV�GY/!�gI����dB�� l��+y������
_���/U{����V�E%�&c��j�B�ަq���ي�p�HCv�]vr��O�s�n�c�_�t��)��D?�8/ �Q�ȃ��j��A�����r���\��2ʘ5 �Ii��}�"�)�a4����s*��e,vi�[+�#n��N�;���Ao�O�ۡ^�dl����'�ϣ����;�?��Ir)l��c�\��¨09XB����&�ƌ�н������e�Lm{Z�[��Z ���U��_C�A�`Hf����m�|3���n�$�2Ro��ք�=��lG?����9��~j�WF�ca������`R�xuJ܉��V�6��L�shB���)���d�Ľ$��ӉD_W?~	.�^�Ok�ңs�es&���Į=���;�a����Nl75!Sލ�Oi6ݨp<�nHhP]Nh�p�?ԁW��X�;��a��Q�Iϯ����Z�n`�����������ξCk�����T&�&Z�c�Zv�}N}h_2���@ȣs{����:��$(F�7��I�����d9R�vQ�)gE@8�]�_W.�+�nB3���Z���C��tb	�u>���-a �\C�Jm�X�C�	�oZ��NOe�3�����2�M�[>y]�A�>HO�Zc�q}mZGښ��bUU�x��%|o4�������=��:���q�+21ŝ.�y�_Q+[�s�t�F���TK銙9���7{N�����~Q?�j�V�3t[��zj�9��䜎NzS�g�z��p��E}jf���*)�+F�p��)*0�����zϩ�����r�1ʿ�$�f�~�<���ħ���������/�?L��gنY���al����q� �2�9|8ح��}\��@������ӭ�ѯ�]O����C�*���_/�ܑ@�%���blIS��[P�~�N^�/��8����dugU��k�`���1L"q�c��4��_�E#o��;Xq?)=��M\<hV	!m����:���ɂ�(y�&��5I~����Ch������I�z}:�$������5n!��YK���*�FJ��8�\��w��נ��"t�y�����
�L�*�l�b��\�[�ZQ�a��v�����,�� io���������[�8a0}�yA��o:��
7aKۏ�L"�7&6��{�q}�(B���O{C1j3���+���g4�fm��e�	Ct��������=PA3x$�����LݖmK��̶��Zn���p!��'�O_(L�a9���@)�����N�Y���U��$;���h��@��&C�>p�Tp�Uڕ�뉲�g��3_�N�BA�Ύm�rta���j�P~]���%.OT�&�:Okh�:���<20�g57���S{���)���Xo���J��e��7�2Bp�w�k[�ݣn?�x!�9Y[�D�f��7M�> m=��M)ތrT�jlN�����u��
�j��x�	J���A��

��h�Sr�I��b�"��
���["�،74,��<AN�� ��z�V��'o,���J��v[�El�9GS�U��{3�����^Ɂ؝a4���j]I)g�)�An�f�{�Y��|��y����2���77@��n�չ��C����Q��a��ˇ��5:Z�
~����S�� eFL`��<ohg���8*]��.���ud��Rb��ZvW��6����O�j��yMm�1�\�P�:p�o�T�T�{��N�p4�D�$t9�te7Hqx�u�uKIp�_�6�ے�OS! ���N�f��\΄��B'|;��r��+!�	�Q{��cU���IǖK�����0ڹ�z�u~�s��o���2�GY�UC��<���<�&��)�9���4��QN��/���/��OYkzk���d���,�hݕ���O�%�7*�~b�_�n<#	�~t�=�@4{�����[P3{knY*SΒ�L��X�ߒn�+S����İ�3J�^�e�M3��|���T]o~�$�MW:򮬍#��|��߃#����$hxj��[��o>�M-N�1�USn���bF��~�xT��uW"�*�\�C��ݳ$JT����oE�x;~����^�Ɍ���u-�
��g,3��-��>/ �|S�5[��f%o�����G�Ά����A�P{S;��ޭY��R�.JP{��M�R��è�V�$V)?U�f(j�ر���W��yq�s���\�:���Y���ּ��~�e9M�`m?���JدN�Ix��5(���c�l#G���G2�ȍ����P	!,yu�5�D��~����u�-AA��^H%�_�c!aR���@2�g,�<�����鿃U�n6���@�槌�gEHD��U�O���
���0k���[���}5�	
� �"��Px5D$w8�Yѝz�C!;_�鲱���+�9��SZgs���X�A�p�/ ���3W8��<0�� n6R���U.��g����k���ӭ��?�S}��ѱ�x�B�T�`��߁L]�/1��OGШ�1O�щ�7�,I�G9�D��=��J=����_��͈�!q(�f�q{`̡�4^�GC�,���x3ɟ�!�l���!u�®�)�=�	xA��6��KM��r�D�ԇN��1x�ߩ�'�)`�g��/�R}�8�ܲ���F����0�n��}�BۻÎ5$��a_���l�)$^�����wFl��aF��G��������d���I����l@�I���?���Z���.z::Rx�Uǩ���g���QS��H���5���c�]?�6��ۦ���(�ʾ��/�6�[��	6��l�{aȰhHL!㉣��9e����'c��Oޣ���F�,O��u*q?z�՜%�ɱ��k�;��
a2��h{m	p~�m���-�����Y�"�6��6��wx�l����M!�׽��g��;PSbR�]�k����}"��|��Q�/>#�蝥�������:T��%�>*������Ɛ�Y��o�T�?�ے|H��ȧ��{q����}��p�޸e�Z]�/btX��Ë?=,ؑ���u��а�q�-�n������m��[�[Q |�H5N?�m�G��]�Y�a���,���]?/���}�FYGgz_�A�8_��| b�[$�"�!ؤ�\��Эr5B��A��Ft!�z�ʩ�Π�/Ú�Y�ow��&�"���T�#^��kV�.t)e�����7�5B�{��9�&
��Ioԋ��JT�q\hN-}���Y�ͩɬ�F��X��v��Y�bĊ[�x�Rϊok�k)��nkT�J���o�~��B mR��`Ǌ?cI3�Pq�J���&.����^�~�{���uV$���1��#yA?��G���R#X��+6oS�(���q�n�fj^P�LW@�'!0N���{z�-VیG�U����������{��BAϩ<r��8�s�-�X%B��W�f����crv[_��؟�����/��?��xcB�e�/��(�1&R�������򭷢D�&K�.���}5�Q�LoI-��,sfF<� �h����G��n�I�[��hpq�� �ࠟ����3}�UOo�gƞ�����E�3�����J����vп'aGVv�����Ǝlz䤲�E�擠�Pw�)����{e��c<��b�M�VLns�L��L\����m[y�L��*23/����@U�'_��Fp�Y}�����G�%����l���L�&גI���v�l/H񀍐��^�:�&qؠ�Q[S#f@x�^�Uj�4ʁB��>�h+&n�ĺ;�<w0-UG~��1R$*��՝�+�oi���ѣJ#�WU���Ltf^������CH�62�?>�<<T�]��t~�5�KBU62��Ff����Iܱ��PUf�|	k�u�F1�a\���>��5���Y����r�	��7xx�����:��*5)��+ߑ�*���os��3����w�ّ"�5=!Z�'$|�YQRC�����}����+�����TJ2�����o31>�!
tRd� �E�=f�i�e����tu�G
�̯�^!���>�N���Fy,���䓈���]Jn
����J�O^��*� ����l�X�ڏ_�S$�@�PR,�<Sᶥ6�6����[K���]��!�=:������{DYG�aRQ�qR�|��OXX)aT�%�䛐E�RIՠso=�ӞF�s�;ع�-v����܏��+����>Q(���od� � ����շ�T��m<�-(�. %š7l�2,ݥ�#��悍b���[�3,�����*pUΐk�K��o���GC��]V�O7\�<g��l��ϋ�ԁ��2���˝����V��+y#*�Xm�xӼ�|���3XI1������V�.�i)_!d��y��c�+�np�Aru���ٽ\���]��,p��w�z��x ��n������S���3B����FC���_D�c���@����O�:�[�l0���+���c�%��ǵ*ߟ���Tu�e>m�<��;�Η3�R=���������I��yG�D��<�9�9���%�ߢJK�c��)�z\Bp�!~�gF6+�T�f3֥J!�^�M�Pצ_rxV�Ȏ�?�{�b:ٌ�5�U8�{�0؇l�
J�eȩp�e����L��,ì�����-NWW�����+�@�i_p�E�IU�@�WX<O���(2!���9�*-S�}ٟ�+ň�0�w{�4C�J�U��	w��NoՀ�CG������L���HC��c+�D��wǺ-� �+�����^�ĭ~-�[h�#�}���'��Hً��xfZugZ������Y���]��o#���%�4H���s��!Q/�@Hj���.N0�������pQ6�x,ڸ2��D�����ME�"?0c&*]
oɏ����n�7�N�%�F�&t����w��/F�I��X12aJ#Lֽ�|X�$���+���
��"V�B�_�&�����J��i�Y��bQ�5J�R)�mӫZҝ�J���cA���k<�<�_�qޒYW��q5�{qȠ~5�i�M6z�����N��B�R7�J��@�s[t��J(������|9��z�5��Z	�	��ᇽ^�}7e�7�2W��nn�O�OK�Og�_�>���-	U�@��&�~ H.Rr�(n@F)�{���ޜCZ����gn'�K�V6�B���f����#�tO�Jv=�֑)�v��"�חG�O��ɝ�t<�qX�Z(c���S�5��F?<io`2`�#Ҋ��L��mj��&[�Iv)��yF�n ш!���
�E� �ú4x*�Yk<8?Yi���82cC	�g�ǂ����ϩ2�?����:��NND��c������6opx�j ,4��._�5v���}���kb��qO�;qBϷj����	K!�N<�R*�g���/��^Û��^6���ɥ��B�e�Z=E�j���:��4k^z9��k���͖�DI�!L�kO�{��������}��罦7�������7�R�!~���P��O;�<(<�O4����6�;o����q�iy������A�
߲2���<��ٶ�-�8����QEY�n���Q��-s1�d��Dr��V����] qN-��JJE:��"d��
��L�O�U�L�a	��w�r~��Q�N�'�U����~<)K��]���J�vRT馄& ���2=E����S��!�����>H]۰�]q
�K��ͳ���� ��D"~-�05��iqZ�nG$�_��װ�L��+�,Lj������Mſ�M�&O�	=9��ٯI��j��!`,!ؘ�t�
��1�� Pw-�"r6��[��Wʗ�M��SGIN�-��F�2�O)w�aSꉣV�λ���u����3���P����F͍W�s�<�l��kKQ�y����&e��/TmR4:b���vxw`D���N�����UzQ:��c����Ր�]�{�z�U�C8����S�o7�~� ��#)��-P�[s�ɝջ��y�f� acɠ;��Q>d�2��'z|7)V?f˕6������e纺�I5ܵ60��[�"���� ��ж>ֱo���1���L,���^0���� �X0Hps�]$ț�1i�G&E!�^�`���*����f�@y�~E}�^�ήO&��b�6�g���U&�,�L��#n�%x�YX���
i0�9']ay�r�ۺ��A{���%~���.�ur�Q����ﶒSb�o�^��3��ޝ'���0}����1�*,i����|�|1�;a�7>|�4��������4��ރ�ķ�d����Au1�C\�,�3���F�T��l�;+eǱkj���OB%�6p�����	�(xt/�׽�E ��0�/ZW<;�g�p�xK���Ӡ��M8�Q�\|��E�# 3p�ٸ���G"'�}L��﯊0d�q�f��,ϘSC[�e��ό�d�T��S�����++0_ih
���Ϛ���|� �JH3���i��A8Y�2����@��M 5��Vt�A�`��8@����Ò������:,Z��H 䃵�Dy���kL�M�mj�فa�Ba��	����+�9_�l�0O$���y;Q�[%�pT�ӬV��(Щu�njE³��b�t�/�M
�(o��0��I{>��i��Ɩ�\�,�H@���rE��cg�iu���s�ac��o����e~;G�#�E��Ԯ��A{ٝ![����>ֱ��~�ҹ�ǒ�-���5�Ҟy</B�ɢC��C	Q���
X�����������c;�Ɔ�+b�B�8��+���t�@�[}/�����?Ə|�#P�S��#7N�P= ����o��
H�2i�:k߳���F��rx�ʾ0{H����>Pz�_�#u��M���C8�[Cw��*���F�i�9��B�5�(�ӵ�7�����ܪaT��Bw��]	fCq���qg_����	������n�M��Y"^ﳡ���z��p8@�n�o���j���)�E^@�W��i,��Hw�X~�E1�Z�*�ͥ輁���Q��ʎr��P7�l5, ����A��W�a�y���$i ;��2g}I҆-�Ks�B�oE�[��c2�="�Lgʪ�0�l�l��Z�LԲeo[o�kU�n�����>e�@Ƃh��޺�~TN���3$��A!֛<��wU,z'|�΍����`
&z���N-Ƌ���������k�J�g���|������~?/��:s2^��+�rM�h_����*7�Z2FR�ۈq����8�ڷ������=J�F��7s0�X�۬�!�73X�x���8��=��=0���S�6�+�gL4�� �Pۄ���,#(�g��!_�P�(�D�����\`m Ԩ.��#yenNMk����|<��J}s|�d�	���_���J��k�F?�
�g�B�J�F�D	���_�Bw�>�*��[F�0r��*�l��$��E|==����Σ^�s]�MU���i��d 2�M)�� �뀜x�О?�,`�N$��P�5J�+c�]���9��-�t��M�4t+T��w�0Ш�P�}�� d��g�����(�*���.�T3�)��q���vh�X	J@���t/_A��]T�eP9����}�x�ʿ��3a�r~v��2��₿�b�n��g���t��`���ݩ����R�w\�s�5`����3DN4'�~���OTzɜ�p�|����=�����
�t���i���}�|�نR2��ES���_�|��F�Txsq=PM�N�p���W���}~cC�f�q�d�|��8�M�92bdl��ܽ���m���H��_k�!�x±be �G�T`���9��1��39E���ؽ2�n+ٔ��C�$�����Ҹ�,Ƒb�j�:� %���oB��v�2x���q����kyPzc��\R8:pا�䇵����<�'CQ��R�ܖ�l�E�#��Rgs��T:�#�
��SlSoR�}�<	7��=��-ঁ� ���(A�>��_����OLp/0d�B4�6ϫ�ly�F+�g��d�؇`�-��"��W5����2�c-�>y_���98�N��y����]T�� �×:���Fs޵�O�c���)p�^J��I���G�����յ0#�ʻ�F=�[A�bY� 5;����5��g2���'ʞ��<�-�����n�Bh��D�(Շ�<ؐ�96�����vT�s����F��.i+�9��9���{'>�憛:ꑩ�a�:�U���/"h��Z7aK����5f�>c�9�#�u5��jA��C��p����I�|�[P�Bh���d�^�Ҍ�|W�_F��2�j�y�N-J�.1"��͟�"��%��d��<�����mrVɧ˅}-ۡ�+�֫�	k����d_�Ѵ��ά���~����ipl�p*D4�ӿ��7f�ٴ����[�K¿pR|v�N�|��1c���.�~[N;~ɑ݉�Z�mPCI��Kf!G2b�^�''��
��\��?���Ns�w��v)T����g���	�����F'�r��V`���鳵v/�Rj�C�alƈ��f���,�W�r��b'E=�H��y��ߑe�ʢ�N!�P�<p~������p'M�F�v��;V͋��v�3a�,l4�ɲ��_	�|R��@:'�Qb�9T��z]P�_O���l(':l?�ě�����	ح����F��!M:1O�h��&� ����5+����?�������/���k��6~��D�Z�Ib�������D����\���W9A�.޿��7�;�{�d]�N�~5�� �F #�3=�.�&_��O�йUG#ϰh���;��f��r�����j?B���z> HHZ
U����c�ѷDi����7������?�/�ӝ)�l�B<��������y��o�9�ͻ+]�����[a֝q����و��]Z}�fPp�}�c�Z��٭*�t�mr���GM�����P�#~>FV���roh��?#z�gH�� �Go���)�����h�SZq|�p��7��E�[��E�������(K�,�<�K�$yPlS��OT���U��)7� �V�F�Z�E6���Ms��PYIX�qJ鶺���~ɍ�%3�"S�%d�A!+�%��U!�b�V���ǽ�9U�_��
�P�ڟ��EFtp����
c	��i,�?�xm����cc���7`�=�9�Cͬ��=���]]\��}"��,�Mk���;u��Ɖe��m�>E�y�S�;��I
Y�<�uw�;�N�Y�;����Q��5ǐ���?n�ɱ��wb�Qg`笜���o~:�X�c�pQ�����^���a���1�Oh�i�Ģ�����u��zMwXD:��*��H��'+��l��<�&>�az2ER4��<=��0TsB�>��W��mq�8+ޑ1-u�(k���#��������1�.#k����R-��/�4��8���t������}(?�'">)��N�)��/��Y�anx�ķx�˾�n���ٔp*۳�d yvp�%���m�����u=<x1��?4:�Y�|���ٶ�/�)y��)�#/�_T��'�@��������70>X<�!�{@?�/F&�����w_>F!�>�]���+��kU~����W85l�2ɥ<��c�ieQ��i�]5��[���?���i�f%�KKt��N"~+��S�i���b��`]��V�B�o	�o*]�=�Լ��R��K��6_���� �{���+�C�|0}�m
zK�KQ�S,���#&�b{򳩰a�Yn����3�J�H��
[z#��:(1}��a�^��G���F}��۴D�,l>/�\Z�u"R�n[�j8��Qߝ�n�h��c�^������р�p����g�J|��k�nM��q!�Njo����=�*���-�{�+�0�"+'?m`�V/1�;V��à7��ly��ؽ�1C\��]��2wJ%�`t�`�rb"_x%+8��)>n�n%o�;�.Z("�T��)�8;b��/��_#|�z�'d�}�OR���%}�C��!PP�����<��~�p��^D�7`�M���y��t����W6U��O�`ݫG#����K�TLĹcS/|lS3|-x���𶵜**[�t�N��}��S��+5>���IZ�� jO��b�Lo��O>X��0����?<��I�H��m�.��T�OΞ"��3i��
BW�y�_��Ã��Z�C[����� O������h�(�(��W��G;#����4-;���^��78��ЩXJ���v���́`��;���2i�pԿ�.��W�n3B}K
�66��v���k(�)�ug��w}#�p6e��/���Q����������2��/��N!�P�	�̓;��-��q����*i��I믏�������"��׬%�N;a�x*�� `��r规CH�$����𽻕��d�"ZB-]��_��T�=3 �Oq�=!�Qx#��&���'_F� �F-�U�{aHC��d��#�.���U	ġY�5���Z�b:]���bE,8�U�RF��	��876�~�ܣx�.�<ֳB�P�m�٢�kX�[*��O��tֻ=V���W�����H��ʰ�:0��*2U��ٶ�J��'�O���3[��cL��6���w]����`���J��'O�.�\��s �ɬ�G�E e�<N��j�h�|jr�̗_��Ȥ��5ap>�������)7�ї8¾sB]�ο}�^�������XWŦ��&�&l����N��V��Y��Yc�A����)�E��+X֜��?m5}cQ���Pr����$Db����D����a�WH�'����D�fM�i�T�F!V3-�PMI�f�7AZO4�A3j���H��U mXR?�ձ��HP~-�l������u�&�>�M�N/8�]�ɪ�������!�ƾnWK�F����׫ty߁"��+��V��R�����%�8}I��Z�Z�e��
���ח�u7#����:;�D�;fU���A/H����qɹ�%��[�@5익�6�z��;9�^Y�E)Sj1UN��K7<���7�D��E/�La5q���w�8̨?�ab�>�/�;!}���Ȁ��%��]3�;�{x����	9�����%5Z�pUiL���+ǔ�5%ɥ�}���ŉ���	���ss��s|���d��*]�����_J����� ��{�>Ӯ�t���H6���&2�u��pV*�UJv��F�V��6(�3%n�B�<�G��~?aRX�|����+�F�gA�>�1Zq!���=����T��R�������Rh��Qp~��уq����B�x-p;��3r��7Va��V�Aߊ���2�D�߄�<}筵X�i���zxvf7�ۧc!}o�
3��"�}�~5��v|��ɻWz>"]CR��~�L��~S�Y�V�� �X��y�mC_���;�ř8�pn-�,���Ie��Kp��VC���s5�����`"JXZ��8V���s�|�t�%�_����7@FUXN���OL�u�t]L`������n�㏒ͣd����DWf�Z<��	�KO��bkZ�n�V�k����^Q��.�#�QBM�q�-��s,!u��n��*-�>
쳑
5��&w.�o�R��pr\㢺@{��1���i���R�ŤK��D]7>^a��3@������W�b{2wՒ+&<(�$�Hnp[@�+Ml�1�[	��\���Ŭ7��e��ʗ �X�.����	��$ts�O6/��!�m2�<���k������ͬ{ �O����V#���/INm���A�eOR����"ݘ�E3����͚�"qҍS��}��=0��i5�9�������s=��۳5ge��H�c�T���W�t����|���ʩ��3S=���|��QPT���CK^��2)#�������X9:����q���v�q��� ~�%�ޣ."��O͗��ٝ~g�RƂ}�D�� �D�\>�O�~��^M=F�Ը~@���Ԝw�<�z�u��h�����=�ّf�{}
������?dYLh[����`l#ʤ�����˻���wU�E����jRY�".�β���O�D8�Rrۿt�qh�8O�������^��C,<�If7�v{˜e�������`]�j~��	a��N�2�ׅo)�m�ۍ޳4��.V�%/�4���?�'}J�A��(�t���gnz���[�q�i��W�l_2BG�r�N)�9���G
��`�'S�su��3�M_��G�?�wo6֏T�~zû��?ws�<�j��˱.r��!�Rʷ������~����)25"x�b��5��m$252�~u@�����1�a�Έ
N!!��W�U�'�_n�3^��Bڻ����g��B��5"E���W���ך���y1F;�V����`� ������3�PBClGkF�G��4��\�x�����)1�ܺLbPӰ�K�e�/�䷱
堢@Zs��(E��j����6%K�_7��5*�&6t2�:��LxV���s���J'�J��|�U�ɧ���	\�
��d>�IFA�ɫZw����}
�N��Ԇ���fG�Y@���pa_����ӓ盍z#����[H���j:RM�y��sb����s�r�m�yUE�uVh�)=
	�Z�͓����@5/�$)�&�,it�oEg|����b]B�8*�ҍϚ~���k��Y0*�|��BSK����n�\-��{(���}5-��?!Nz�݋�ƙ=$���,��Ơ��3�Dx������=�%�6"��ƺ!�b����c`i��2ŷ*\��û1M�vtM����b��{�)U/1Qӧ�Wt��ִ�K���f��O�s���=r�
�P93fK�+%Hh�YJ���N�Oz�?�z�,mV�1���5г�����0����^��q�k�����fy�cp�<gD��1���iʩqDo��+�b@~ug����Su��ȘC�E�s�a��ϝ��.��������b ����籁��WK��u:{�-���CvE��9*�g�[ޑ�D}�ڋ�B�)T9q;NHfb� !��e�&Ꮬ[�%���w4�}�}��a���C��{"g5����5I��~�L+S�YRf�l�Wi赞�$x�P����#�r�ԁ�D&���Ix��ֈR3D��Tп�ʹ��X�s<�5�����5���}�x������P�7q$�+A�#o���d����N��&�$!z� V�����3����ԁ� �����Ŵ΋~,U�S�sy�@*:����,�`�v����ѧȞ(�S{81^��p���o�ã����q��j��ݭ��63a*����N�:[Gi(C�xŭ�ʼ[p��/��My��$����N�{��u|5��/d���"��ԕu%#U���;�%z����]�vm�)C+Y���S����*>��{�2��D0�y��;�_��s��'�����
��r hs���=6.�p��� �A�����U��N^z*>��;m��X�А��N��E����ɤ�?٘c���?z��k�=lݏ�s��֡Ĉ�IUwJ���F6��J՞܏�����W��f�������e�B-�F����О�|��)���?Jt@�.iSΈ�D�V9.@�BS�a����۪��'p���OQ��Zy`] �u�͎n��G�=g��HM/ATq$���;��a_�>�w�P��<�c���u�͘C�m"x����*�*C��E0��Y�8��q��d����:����Z�!���ZEh��e��� * e)��g���^��o�T^���g���LC$Us��X��X��|��g�w�,2�T���^�vo��y.�~v��})$�}J�?�����^ŎGE<R��C�y[i6C+?֔�]�x���C�}�Ķ�RV��m�s�����)G� O1[s�L\n���g�QK���������F�;� �A+5��G�9���͞;����k��� �v�gV�C���ﴫ��*JF�p�WҺU�.K�)S�rޠ �)�]H�����Ş}2]	x�K�]�V�΋���+����߁�ęE���ێȜ�þ�+���S9R[,!'S-f�G0�����%(�Lhqa����u/B�	jM�8eq�q	�fR�@�U�cZ�q���!���l;����V�{X�P��h)�jӠS�pIBGm=�?��F���t"nn8`,�4R��"c���Zhn�Lr7��b���ؾQ8�T툼����!�`G��`vx�6R@��:�ɝ������6y2��m�%R$ʕ?뇩6��~��j7�	O|�h�I�͹hz�	^wF�С�N�+��sM(���W#��,���J��
�7�8�����[Ѹ9�z�L,X=�+���q8,Qc�vng�~r\��W�~���\ȣ��]����V����s�\���?L�����(
�ˀ����MQ��.�S5v(���d���4����(W]�/O�a��<�~dԪ�p��S�v�g��fꡮ�H�	��Z_�շ4vH��g#���Gks9�(U{r7��< �*��R�������T�Y��,H:o4[kn`$��C\"s2�R��{��pQ�9�����2Z����lA��G�=墹U��К��@'�,������1�-����tk�Е����M�����E*3�Oڪ�5P�)�'���;kC��d�@��\��m$FL��xY%�d�ٕ�ӆ��V����Ў3X �3n,�͋(�+�GqC�bï3��Bg��R���c���3�~+�.rθ�zе��.-�z�ٓ�ӣd�q���dD���/��9���8%_r%w������O�=
ۛ�4?g�8P`�Wa�z6y_�#�a�,��VQ�t���<�'�����=��K+�k^��k*%�/���>�� �W��:N��.�	1�m��<�c��8�-�8�i�z�2;�c�'��3�eI��#�� �<��+�M�$�neVdt��Y�b�
�	�rj������ΐ?�郵��pu�X�z>O���y�MR�ɍ�&'� �\? 6���m?�+p$���^T�2?���O�m�l���u�������b�]E?���j���j��A�ĕ�$�Ó�&Ηk�y�����їj���fa�:f�/3֖p���'!HQ���Cj���z�!+�1�۫?w���ҶXX���%���T�!�d!Ɗ��W���gqxVEq�W��m�E^7%v��x���qf��P2S�������=���Z/��<�-HI5wD�-d��"6 �q���my6e0%g9��e+��/_\�DL��Y'�������ޚE��L�$3��'4�����mY	��z�Ҳ�bftj��I�lXL79�e�����ǹ�8�O"�imQ���+(��(S��=���1g����&Ò��������O:Ϯ�u\����^�Ѹ�T�
J�+[Rj��m�C�"�@��Xe���T�ﲍr��F���;Z�j����onn���eq�C��i�y���Zě2*�ND��옌�OD�y�˞��f)	ի���V��V{���?���}
0���v ��Q��R�@X����f>���h>�\��,A�Cw��q����,OZ�X�����]z�ul�fҐ�Rz/+�N��XcZ��u�>���6޽$K�̫�M���0�\�72QΞx�c���d^��{��;�6�ϟ,������eЭ�{����HF�3�|��L�kA��������D��'��&)H��������E!ߟ�'5������!�i�J�V�fL�"�t�zՐ�pk��N_˰׹t����)��@6�)�{X�ǭ��W_>!L�ɓB0�Z��������^�>Md��__��|M*��J7p�I3���}��x�N ~HS0挏�,[�$w����0P�M0�i��/�1��iw��چ[k�� �ui|�HY߹AY��Xw����>|�iG���|g{|A�ʄ4=^G83��ca�f �	��F���%$����ac����7J�����Ulс�W��]�\ޡao��/>��s�NW�>U��]#���cY| ��\J��2Z��O��쟟-�����oEQ9��N�l���1�+6Y������VE	[l�m\����J�r�w�-�6Z����T;i7L#bV��`a	
+G����Y6ީ���JfZ@�}����s��t�<���X\Gg���}V �TC�b��Jc&�������7�yv��凞�W�L�S���xY�9��q�û�!�L����A�i����P,�'z�ǹ"6�]�&\M���;*j����E�dj�����P���SÓ�p�XS͚2�c��
XDҬL)3o^��9�Ț�;�u*�I!C����&f���<C����on^mB@#���T���� C?��9&3H�	+���)6�T�i娦Ћ���8}�V�F<?r�1�������į]{�N1o��~e���&�Nt��1�"q�냐ͦ�d| ��B>����ƆS�]}J	��*h��	�A�Q6/27%K��u�x��7i�W}W���._PM��繨���y[��>��<��'���t�.�0�y8?�Lo�9�p�Z���ӌ��/'�m�(���'�J˽���[���>\v�Z.^LX��~��-Y�J'�w�ѓ5K�� hO���}�p�"���.W}^Q�ʮg����	1�W���H��|�0([)��s��7�j���*o��((ߣ^*-�$v��S��6��f�"����y�����M9���}K[l��x"�H@Y�9I&�4����0�=��p��m�Tx\��Z�AH��ز��?�y$��ҳ]��W�E���0��]�_�{d�N�"���'�}u�aNp�����A���'����X��&1��r�;^x�HF�{R���u��p�(��OK]�4~�Zݾ�/��۩�8��C�}�nu���L�0O$k�3��b>Z0O���U�{FX;�sИLIۑ$=�ZF�h ��m(\�Y�~���A8��������w��WY���i�ϒBkșF��d��ww�>Q��ޯ j�^8�x[Dڮok`n�����-�`�@�]��W����O����h�L~\4(.�}5���gP�{)X����d:M����H��HƳ��s���\ؔQT����1�j�]�$P:T��m���Z��3��T<�o�Lů�W��+��c��o4b}ЭD�9Dd�R�㉋-~[���e�Φ<���Z����.��Y}���
 ���3��8Uc�vk�����|_�!UD������ҖQ��<<L����Kv^��	����?0a7�!5c�"�J�y%��ȱ2\�D��E���V';��)��kX��n�n�d2a��w�u3	V��9�N0+���:��
ݭ�j��e�%u�'�q��<r�P~�]/X�j�f�O�/�G!�J�T�P��E,v����k��ˮ�JBv�����;έ>BN`.̯�7�@�/|M�x�u]��W����>|���S����р"�v9.Ut�ε>�T�:"�bѹ�x a�DC���:mҎlF���֭���Z�)�v��ea��ow%��Ģ���ZƖ�0G�_��Z-Ÿz�h��+_c1,�(̞��>G�L�>%q���x�+����&��6�:o^k,�]_<u�cwp�v��J\ �3v� �=���J�2�1)zhӒ��CGKҁB��I�p1s���ڃ7|�=��&`K�⏆!.r_��j�>�FಈWJp��$?j`���&8�j�%��	l�����W�8�4}��N�G��X����G״��ebzJ����u7
�,�C�/�(nG> ���D� z�WD���ݽq�+���@��{���Ku��4R�g��ǐ%��u��t`�[E�D��K�
�lsY2�n��a��	�Q�\��q�8ds� ��h�V;d,��w�8?�!��"B	�>_��)�`�:Z�"L�7_$Nc�dA��戃�ӆ&���-3M���KR~II�!7���["�d���	Eԟ�e��O�"���H�q�����rֳ�<B��>�v878nr�(��q�d�z!ƷU#T��άۆ�QѴ��ܘ�cAp�E� �,�(����☱.U�Y׮�N�P}̭Z���(�4��{��L�ʅ��OhF�.��;�����1x?G�t�x�ɶ�+��99o@��7�Ȥ5E'�����D} m��BJ�A��7���a�Q��G�����.��K�O��C��pn�]|EviA:��9Ot۝���_�����������?^��`�׾�%fc_C����3BYG�X��F��,�*I���ɒ}f�ʖTa�R�AK�|�ݿ��<�y�߯��}�9��8������h�>����H�#��ړG<s��NB���r����v�6a�nʿ�G��p��<�+ÿŞ����d
������]��������=G�[*��>�f�<+����nQ�gfsE��T�ՆG]W�.3�o�
~eK��2Y{c���d�Y.-��j%���nK��5&}gT�Zl��d���<����O|P��!���<{x�/A'b�v��\��!6eP�X5ϸ���.�����?��\�A�Z��̋{�Z�����[0@Xk�LU��X�i���m��kK7.�(���X���աl�?^��}yn!K[4V9_�R6�m��iеp�1�lv��Ͽ|{I�͏,'(ጙw�g�ֿc�J8��S�q��W��F��K�Z�)ʤؿ�:�Mn��\�U�;�U
bF�~R���3���8\emH�g��u�'/2�^�<�0�G�	;�g(�¥���^I�L����_��LKҩ��c�<ҝ�a5�nUy�2d��'�&-y"��e~}�?����D��(v��z2�
���!ּ�̨��ޒ"joob|�)a
���x���� �3%�Vi�M��U�lu���s�hBt�کb)���C�3��!_4o�+� ��S
3�b�꥔�Z\W��p�Ʒ�8�z��
7'ޥs-��{����C}��í�z�S��p��8�4�}�T��Kl"�zƫ׺�Y�m�GjY�����P=å��^=�����kXIn�4H��%���wڢn\��i�w���Z�-����2���!�NfZ�=�cnk������Ǯ�'�z<gM����~~F<a�:��v8�4Sڗ4-]��=�t��yr�}7ix���7=���W9�� ���}�C8ТD\8$��=��=gU~�@�Ս�K���2Rw�嶈��!�p$>)S�Щ��.��\�wQ�~ �ڎ���@+�д�,Ę�JZ�/h�M��)�_�̭_:#�"�W��]���w?Ol�2B�|�͡�<�p G��A��A_?i��H�'�[�C�[d���_�789�( �=uϖ�B�Ca�w�T�G��
\Y���͖���s��x%��{����<�gvڙW8Y��b�іAE��C"�.]�t��]�k�<W0����m4j5|Z�6�����ďn5��I#��AL{�?�ɵgF6/���~G���"��W�l��I�bs� �@ג�ҥ=_LJYA��Z=�������T%I�p��ö�(�v�Hߌ����	���\��~`\/[0��^^���F���%�xek��j���g+�Ѿ��Zo���F&�Z���+��!��Ӌ��+ņ��)a�DއFC���G*�W
��#CS���r���Fl��ԫm�]b��*_��օѼN�N�>��{��»��!�����H��F�d��u�F�k�[����������(�x�L���9rN+ґ��&��8�A�G�c��qhYg���?���b秴�Ty���-ڥ���yj"�k���z;��m��b{�8ikd�zG�Y�)�F����	7�Ŧ�B���+.뼑fq�Ѽ�z+��^�N��H���z^������ڐ)����r�(de�p�%ނu/x�/ܺ!�q����W�R�AI02Zj�ls��mp�5�J�E���D{ Bu ���;���"�և�~�נ��}�W����$��r�X0H���>��*�s��~F|v�2>A���LW�y���+�NLH"ʠ�	q�ZH>�MgGʸ����w���ǒ��LO���pko����cǏ��v�1�d�g�}�����m�Ʌ���Y�,M��ii�o=)u.�`6�ޑ�`��Tfq�����C��m�����W��x)�����#�CQ�Tr�[�%�<�����h�s�B�ٖD�[%�#����WO�n�����Ӱ�5�o��TDX���%���lږ���R�=Qw�����X2����C�-}kZ�Gi��z�@�?�ݸNN�b��J*$��l��I��$6��w�w-r�[��_�������6��.D1�=��t���Tw�3NeI+��F�e�ƭ����n�,\�I=/,lj�>��V`��g~�_�ٞ2��6�ÆP��z�#U]+��ܑB�@N|�"��7�m-W��	��<8�R*��m�W(�ޟ�;���T��'x7���8�M;���P�"��i{X����x�yF�1Su�o��!����R1lӱG6Qq��o2��*P~&�|�����T8t���w��Ù�2g^��7L��dXz�B���,dx(��Tlv�kq�1�x-��'�`1e��ـ���|�8����c�.�$2%]?���GZo?"�JkB�x|��!3hܹO��GF��E��W�J�KW�wk���]a=��`n��_�e&WÌ�sЁ�� �wn����	Ň��J���8y ]w����#�RRcR�M���R���_x�!�pU-Xh: �t"�V�(�&���iIiZ�����&m�����볮���U}��`�X($��,�ح�����'X�������{�^oץ�鍶��&=��ֵ��"n.�RMq��U�s�v�PBնK��?����Z���a(&���ko �z���F�s�ͷ�=����f�����E�[��3����!���F��O�۫��/ral�����ɮ�	�ѱ����ȫ(�f~�v8�����00a}�Z��ȑ��u
�Ǖ��z'����}�v�?�8롞��VJ�kZJ��U�"x>��薁JFv�Ɠ�Ġ��X���DV ~��Q���Ɩ_:�-��5�k��:þ��0y�)	�ҟ^H4xC�������F�L0���>;p�����c�����s��q�|�)$�F3��[el�K5Zx������6�}���z�FȒ¶�+t.�V�3Y��Zdj��\.BH��@�ؒ{�MN�3���0h��A�L%��db��x^ζ2��U�w�)��q4 S�A<�0	͞�FLMC�����h{��L����d��2�ʉ�W
n޿d�O�M�H���(���"��F^�L����㫷M�y�TMi#��4�6;R���6z	,�}M#gN��RQ#^s[Q3>4�:������.&A��e�[7�U��q���ȧ�W"���$��[���c�������nDo��x����h�勖�F��DªԺ��ɘ�,�#b?��z�kg����H<IuW�$�K^Y���W7˵����9#�S�"�pu�R�������\�9�_g��^���~�r/&����	�kͬ?��+�>i��v��un�s)��{�H=u�G�/>N��ы�$�0�7|O����.�E��y��V�\'�^�h2�����z����P��d�-+aXWGӒ��w��+�]MlDt\CъJ�����������fs�u�2O��U���Qd�cR������I]���0^\3�Zo�'.�K�=P:�D*�G�L�%��������g�,�mh��sP�s�͑3�mmf����
�.�h�����C;``���qJ��i^%��-]nK��&��NK3��=4�b�7���`)	��È?q��)ﷴq`��z/���0�$^1���vm���.73Rvm���a�O�ԃ�S��-�Iw9���CG}�	��t*�j���3(װ�s�p���ܓKP�C]��Lsyo��R/�P��%T��<0b�\2�/P�Nxޯs��p�
�^�4Kg�_��\ٰ�c�*FQo��F�LMP�>9���+��[*'��z�an�>~�$�y�}�z��C\+��:�_���|U}���%������J�:ib�� �$�L�:���J�n(�ڙ��V�Jƛ�����=F�q]�-s�]�����c�R�¡-��l'�,$���L�'�����p��]0ϴm�U	`]��>�����ѣ_��s��y�L�+x�tJ��������2�w8t`�c_o8�i�,b�T=���ٻ�mq������#��ԆϬI�{�1�|Z8���24r���:�J,��X�#��a._Z���~;���������|OK3~��(cȄM�u7�8_�����<s��+z�u#g��&�)!�FT��W$���Dh&n����曟Wwgc6����^���V·���6+���vl�ON�]��;�3�34���/%~ۋz�ȵZ��xM]�K��i1����4��n�b��'`-d|��G��fPK媟:1\¯=\�ݖ-h����L(<���n^^��`rn*r�2���'J��~�i��LLb�H���{��#��[�<+A����Q��H9M1�o��$�گ.->pD��sX���vVR�?M�d�0x���r�eG����1l�sk�J��NnB[W�	n�����~B�U�|����6�@o̱���	����S�ňҕՏ�ͷ8I��W�*��S,�bE��v3s�ʁ�E�أ�d���Re{ECj���pq2��PCD�a�_���y�4�͈�҇��T����7ι^�cT˥I��k�j:�ufx�4�v:��\-_8�/�{�	����~Its�D�U�9���O���ߙ��!D�Ɓ+m���4�2����&�3�ʗz�'s}(O��ރ���$6m8�y����Ӡ��B/�
�m|f,��`ޒ=���y�ˠ�;��=�6����-���~=5���n����f_���W.���:�e��j�\�^���68�����t9sVp�%��V-�u �s.�&d\��5�g�:I�UhP�H@W��Z�RFǴ`�j�E�i(m������2d�~��U�j��buVSX���W�����m�e����v�P����x���g�|���v�s��[t����"�ۺ�]�x~�ܿF+�l�Bƙ����KŶ2#i�=B�ec��2�&V_X�(�@Tіe�7;s�Ң�E������H��q�dT8l`�p�z���^�%A_��\L��s�-1�d�������)��Q�\�܆nN����مbD6�Fr��8zd�b>[k��$4�80P�<����o����XB\��m+9)�5���2r߯W���cq~��sb����&p��fa,'��u�ڋҹ�N������#�͙�i��N�3���3O|FS�����M��goP�EY,�-�]�a]:w�[�[4C{w���]g.���ft�:+���Q��3�\�r�/P/��ʶ_Z�1��	��D�3tM
*�
��
5ˀr����kV%��4
b�x%��S3�l\�1�vE�����Jl���V�]����C���f�@tE�+�Z��4��Ixe>��2P���@}?:
_᪸�<:���}�a�+>��%�ʦ�*�H����:v20����Y�uj,�`0w	�Ow_���߷K=��
S�Q�����\�j"�x͔��yASo��vU�vr�~�T"Z����1�[����5��\�O5EF�)�#��Na�5noz}��,���a��ݚ
,k�bḪO�*%j@x^Ծp!7
�َ�@'�nK�V 1���?���D}�U�����t��	�Fq�C^ޔX�u���Jj@8��K��]y�=�;ߊYT����2�ò�#�� ��C �k:����I?UuXC��~��î�z�YdwV+ʸ�V��z���;��.������H�[�,Ud��6��&+�̕��_�5�m4FFJ�g�U �����@����X���]$¹Jg.A� ��hӬ cW�-���f/Fk�7�����R0���zw�x�՛ǉ��p�棫��=j�\r�ڋ��S���4���
&SNk���XJE
��}g��31��R4������?�J�d�*�'p^�P�lO#H�ۚ<�3z��	�vQ�6�C1�SKe�D��"�r�6����JR�a{�����]�O�7O)�������4tRT�^�����y$<��P�G�㳮79�����,�C����SM
��S��n��U�˕d��34���Yk�A�!�Ƅ�ηg�c����-�zm_�WK��L)Q��MO�o�:������y���Q�X�}ZLV�]r��P���&������X�2}6'��7���UD3j��pv�	�Z���Qz�a��*w�=v��f���S_u���]���c�
��]Qڟ��"�דh��%��$fD�����cE�>(���ڽ�҅Ċ�/�;�ELdMV@c��/'�r�fK�ݏ�X�s����G�D��La��6s��p�k�%��`�o� )<^�9·3��jCRq���gao�����^]i���GܠH!�r ��

+<��ӕە��U�2�~К�T�QSeq=��z�b��T������^>E�k���n��V��t����*��T������dO9W�����S�Etơ���a�)(?������G2U<�͠��7χ�/uӁ�>�\A �s��2�r��{$��I;��J���?iG��0��"n6�C�lw"m����B/_�خ�uI�j��h��V�8���}n#���)�d�T%�(锤3�;�R\sw��%��P�.��U;L<z����4ݣ��o�;'���Uh����/-uK���_��)���Z���=���Fٴ�ԝ���Nn0�����Ɏ�>�9�DjOx����A`��Xi�K)���>�����p�3�a���%m(O�(Ske���	�+QF�m�t�w�c����pCKRNE�/�W.��9Һ$g��<ˣ�?���ƫFP7&~��3��<�ǃ��t�;�4�:�o�
"J/Ax�}�Kf�=�XKA��%T@YƤ=�ｕ���"hd[zd}���X�׋��C�Ac���q����x[m���?��i~[�/�y2�Ba�C��m�^���i�>�)WPk�R�y����?n8�J�̄�E��a��_t�V�qA���b��;s�"G�+Ӹƃ�'����i1z;ﯻ�E0v0lt��O�>2[���^w���#�6�s
=��T�z��l��:�e�,k� ¼9��D�/�u�ď���y�䘘X���`�I�'n$#��#�<{��r{Y[�c~3U�s-�c~��{?e�W�1�#�V��� �9]��l8bA~���ȶ�6��+￷��(|PP&WA�-�n[�6�����Q?:)�#˗�t�*2��L�+��:4T�ġ��c=v�@J�	�����\ŭvkw�mF A$�;Q1��~m����[`�"�����8�o���������ҳ��*h�j����q�l��9�p(�n��jdU���q��tv�� |�#���e}�:oꉵv_(��E��+�F�@�����X�zԡ\�~��V ?|[��A���	�QOvbU�[��'�!��k�
�0��<�d��V���+��G�S��Hzg���ݏ`�Ho�pm���fV�$76v�q����)�� �Ԯ %�BK�w�O�ܭ%��Wֲ�+�������i��ϙ
OFB�9�F�|8z�>x���hxW^0�R�1��U{'�ӳb:ގ����l�I㉡9{;��Ŷ��To�����+����7�����:zerv?�=�\�H�W��r�������ͣ�_7����֞���ٳA��&~ �[x��`8D6y7w���{��L\R�v�-�`~]^�3aa�B�Ŕ��su}ų�%�"�į2�%Oh7���5�RFBd�W���ֻ�l74湗f?����=H�I�d�D�|��J�e�S �y��i���2�/�[����h���IHi�όO��R�	,��"iduQ�n������Y("5���
��>������ET�<c�>��QL�����eF�>E���q2��[�#��{o-Cg����S� fE�pzi.?�Խ?��%i��
2N|2޿a���������L�w����j����k����l.�\��g!H�y#�9�x��ے[f!�}�M�+)�����b�zsy��Ҙ+�8�UR�0��<��|��ѵ��q��mP��ZQJ�}�/^^%^���鯹ޔ{�y�' ��2ȋ=i�j�x�;|�_+�G�倫Q�#��<�x��*��vR8��w��3����<6x�����}�9�!�i?��� bA���dS&�A�R�]׷�, �8�~���n�n҉���Ϻ���WP�{.�-'���h��L����Y;8�Q�F�h�F|M�B�(Q͡}���ެp܍m�r��#� 
�K��ޣ���P2�uAil1"f�j_%�TE��	;���͊S�����D�yT+��/��P��s�n�s"�Ij�:��>�4O�e��ǟs��w�~�� �� ��iS
]E�djO���;�[������~�r'��S���;�ˏe\ROʫ󙀸6�4}�*����\^Z�t�0��k�h��� ܽB������y�A�5��+�<�M�(.��Nt�I�����
PM��4���+��Zt��1��B����L��3�kP�^cv&}?zgD�3�|X�ЍP�
���0���4J��g�T��ɡ_3n;I�ͭObf��M��j[\���Ȣ�-�"��� dm�ǯ��{*^��z!�u������ާ6�NR���X�T��ǅOR���l�	�D�p(O��ﮉv�v�F\���%����ϗ�;\֙�x�W��ecW�B��D"�B�~��:��(�Gq�am1�>�;��z�2~?�g���)؅475Q�7�Y�'��`�I�\icF�=~�]j�jgH�vP�8|Tz:�ޟ��rũC�����_�[z�-����	#��>��j�ħ�^g����-��h�CgJ�PѮ�|=0�{�0u�7�����d�g�ޢ�{0qYj�=�C蒛����BG�r5<o�Mթ�kP\M�8��������¹U���,��m�G�b9������ *�q��/�h��3����s��p���(���s�+b��e�Pf�#�ޒ����\^u9�����.�KI���4A
u%I2�O饠�����9t��,A� �RiuLn
�a�Q�-_�vU�����,�k���^9��
���y�/o�m|3��(+�/-��Jv��w�){�SQ�:Pa�
gHW�:��x4�����c	�J�g��W�0?��ыY���f	5�㹘M�E���W��~��ҥ�G*�G8��y/��,r\yk'f�-l�����)	/t)Yb]���{W�d]��}D���� ~�N����~OދJ�W�Y.�5{�Tqj��R�2���(��6���Ych�D<#��EQ!.*lD���*���-8�.b�X��A(?��VgU��d(���X�HIV�c��w�#��H�0�H��n^�m	�I����"1�˿"Hv���+qa>ⶬ��j�$�ᑙ.-�2�Á�ᾰZg�3N_��g}��#<]t�I�k��,D�-� 7�����l�?�/t�|���4��K���!3�y��6���¿#�ė,ɲr��|�)�@K���<J�y��)�~���f����uk�fr��k�T.*C�Ѣ��ܨ�G��EL�r�����yF���\
���<F��{#_��v�\��?��op����@�N�d$j��i����v5<f1�?Y�xΑv��ص�N/�q�Y�6���U���m4�������Ŷ��!<8	Ea_�J����M���_��Հ����<�VV�D���|T�,����18�%-C��Y]�h1��;��� ��L|� ���H�sg�S�g�ԭ]r�ճ�c���i�`�� S&Vx��1+�z�j>��S��5�5o�
����kË,Ѳ��a##�Eso�ʪ�o��b(�#���6&�!U�8в��/K�)�G�;g�މ�`D�#5�7-aJ�?V2��(&��~�Y�Q�z4K#1m�R>���իt��K���y�UHۼ���6������+�-�4��u��	��R�+��᪁��Xb��)s��a�@���n5?O%����S)"���؝[���������Zv�Pʘ��i7���W�����|'��M��3M�=��m���.ى��(��d+���� �I軫�(Iq�]�ti��/����B�5�؅�%|�W֩v��~Q�=�pJ�<b��SБ��Q^�ԉ��K���K�i|���Y$7I�7pW\FF���C���c�[��1�d�)�}��!�8�Y7JBC��܀i�$|��dc�;ʇOˋq8F�-m
�YWXf�s&�U2�!���] � U�.�|�y3{���]�_������}��-_�h���\����̨�jT�m�d
��ɭn]]b���ѽ.��D�H�W�׻�d�+�w �l�4��wa�QW\3�R,'�Gq%m��R��uR�s{�8�<9���m^sgCN��ǰ�LN�j<(��6ư����!r�Et\%>9�0r�O�G+vѴy��c���lo��wg*l�\j��ܣ�P�%/ɖ8n��4��"�enKx� ��ίK����hgA��r/�]6ʹ����� ���A�}�V��Z��	�9
w��ř�4���@�l|L�!]לgt2��4�^=Ͱ��	��d'Q�b���rթ��'3��ޕ;SrQ�P�O�t���p(.߸�>���q���ц�AX�1�\�Ȼ���,#z�cu1�	��V��Hj����5FJ~u`zI�V����M��V��:�b��pߘ��!�1V����"��M��%��J��ϧ�棨��z���FS�-c�AG�4�[�v��;�al5���t� �%Q�G������H�ɔ��	���o8|�W���H�q�
b��*5���v�sqŔ��ck����p�4iq?�ed��z�X�2�P�S��=�֥�v/�̵���[�%��`	\
 ���.�HcZ���aP-BYu��|K>d���¦�Sh� B�����0V��˖���z�N�b|�? ����3��>8=a:��4��'�DJ�����Y��ҩ�'Z�I@Ϋ|�(�������^�K�����6h���y࿓�[@y^h��CGR��� _إ��VW��n�/��٧8�*_���?f��6���be�\.�Q��߅�!P[" >�a�~#�zP)���n�'+8��oګ��.Méb�9��wC��?��l����:�!N�PVU<W���R?~ݝlB�i>�����3��L9�jg�ߞyZX��++ӡ?�ۙ��>{�B����?��Qf�}�ɱ3����`�Q����hO3S_>� �4��aa�+C�ۣ��he�(/S�H����Qn�<���U�uB��؟�[`˰z�ʶkqÝW
�C�� !�ӎ�͜�#5a�kx���KVn
 ��nM��%�>\+6?�&����ׂ^{�<���W��Wu�h����}���".B>��9X��>�9Y�OYA�`ĵ���$*�5�u!Ċ�M��"��Er0�bOL���vb�}U<�
)�t�g��`O���ߍ3#�;'������{�q�4Eh\9"@�v��$!��+X���� 9;�to���l]��|]g�fOJ ��1�ů	�͕��.6��dLV��#u��eL�潎�^#��{��O��m��2`� <��5��n={�4�����NV�2��A#ىzNަo����g�l
����A��eE�@	=A+�rt��=�Ӝ����g��nn��	� P��~ObW�c���o
��ݥ,?�AF9�܏�S�R����d����Ǐ���s�ϯ�Hآ�b��A���H<+}/_�1�[�I�s,2R�����_^�����`J��6���9��U���(�3h���Uc%s�V�TCL����1�y+K(d!0MF�e����sc=	7�փw?Y����f����U_�T�ρz@Ϣ k���fTe�������b]3���]��Е��.�)<�,~,*��3��h�5��Y����{��!�ۿ�\��2(Q3٣�h�֪�O�9�TU���ޡ!z�SG����ͳ$L9Q�����8M�%%(37(2^�*g�"���1���r'q�-�Nj�jk���]+|v��#J/B��Kp�z��˒y����9���������\��(�CR)�$'�b��C��b�2 Dd�t�6*�^C�^~{�O�������4,����pUwL^�E.�f�,�Auy�v�%�җ3���ߊqo������#ߑ�og��5��"�L�՛���)��n�U*�Ē���10���+���+�MRʦ�39�} �o�Y�����k?z�G�z2��_�����|Vo{Kɵ�ֱ3����KO0�
��B��sͿ�^���I?e�λ��<eN�-^�3�M4���l��!+��+� 9;�`���hm��-Ge�����:���؃�E#a�g7��l�wo2�>LF����|�hꪶJ��{~�Ӎ3��R�E|qp��pJ{y�In0�^|��Ņ`�D�9���f������	n;P�d�q�(xpq�moғ;�����-?�Z��e�3����s�Y1�]�-m��{�� �H�T�����߶�M�ט�j+���7nU���{5c/P����lʓ�K��j\�!N���*�LDk��:d���DT=�uu7ggE�����ڰ@��fEQf���5k���� ���IHl2��q��Slz8�`
9�=�;��C���_o}U�xfO�a8���z2P�o��=�)�,fas��G@�O�1*}���Xk�*Q�h����b�����f]�C�1ه&�(��wݚk�K?�� �w�X-n�X�C ���G�KE>XLq*�kR�;_�mZ�H�>:�Z�P�ЮV�ăKwT_Nb��\��Q
�u��$�O�~�~\|�;?}�
ys2��Ś��_+){+.,?X	3���^$�x����/��r�BY� .b��9�P�p�c��\�$�~�J%���}�����'�S�����Q��9��ί��PI�8����M��z8s̼T�x�3���Xzq����UM)�4ee>�h����F	)�M���@��V�r��~��N�C�7u=^��G��
�#yj�,�x�^|o*�S�	A���gG�j�͛XCJE�<�-��.D�C(�N�h��T�����}}yz���w9�4��Xz�Yr\��u�wc���M�"��|!I��Ϲ;/�S���*γ��j��=U�ƫ�釵_��Ӫ�\�@�7Īrg�S��A;�?��ն�U��⒤���bk���ɧ+�Y�������Q�%�y�#����h�K�B#\�5�F>>����	�gE:7c�Y:7{��B�b�҉#�,��*�q���>�����\�ˌ����}J���XM��&��*I���f�wu	ϣ>i�50b����P)�1�(��8��>i'��֐P.�2���D�iSY�����F�~[�K�w���l.'���J�9) -��Y�J�s�5ΙO�	����w�UW���Zi�ܸt����~;kڣ��q�`0��'���c+���M�_�{F�����-�T��W����D��X'�Eh/F`�0w��P/:Q��Jo�T�(K���eXz݀i�ل9��90����J�2���UyU�n,�CߙX��	$�������e��O	K���-Q,�:3��������8E���b	+��J~�dx�-��v7�?_��������#t�qGY��r�q(�b�-b*Q�_����_�?^%�����c�����F���D��EX����`�G���OF�"��w'IE±o�h8qp�Cy�Z������ےid�E\4�����BC�Ӿ@]lMA.b�>�n�����kz�N��E�6�t�<�B|pYE?^��תE[�W�Z(BG�o��k��VZ�:�2���M���$Q�������A�?r�� �����n֢�oD�т�aE�\��k��đ����-$x^�G(uHZ�gƳ��o_�����R%�D�KC�HL�ۦ�4��E��⢥��bϑK��������o����J�Aɀ��b�]���ȥ.+�a,��*d�5g�����������-����Ǎ'�	ޫE�7����z&��D�+δ�b{&�==�?��I�poSh���r�إ�H�ě|f���蟩�������Eɋ�&3uvz�i%���C�>�Q�9�=_�W�,ZXd5��������f��/��,]o0�Aq$Q�ݽ���7h�9�Ӻ��Ԥ��)�^pe@���F�fG��l�t������/�QKY�I�#������n%C��!��b���KJ��~~���o5E�����Y��7���3���qv$�A�c�w�	?�;ϵ�#�,YK��%�z�!‣}�)��ʏ�q>����!�>���\$���\"b��.ZZl,��ӊZn0.�Ċ/�reT����-N���֣{��k�$�� i<@V=84�x��ș�[�zsb;�T9�������x��y�V�u��q���8��g�����s��*��E����|��T3�W{�:ܐnU�H�����KO�u����b���TV�jt3��^(��d�"5�t���@�5����Q1[���3;^x�7�[���<(>�C�B�7�־NGps#	���;�����sqb'���j��}O{S$�<e���$1�H ���]��T�/Z"O��Av}�*�~��ɝ;'f�{	���q�%*���g_[�0f(�2ͅ�0��ȼ�����9f�b�O M�B*��wY���o���( �|��/j�>&&a� �j�d�M���i0C[���R���دj~c���ť��τ��2�{����Q��(Q"���ybU�nm��� <׿�Rl^/�l���T\�l.Ʊf,�fe�O�N�.[ԉ>_��.����Z�usDDp�ii�'kXŲ,hd�8��F�U ܵk�_z/�1w~��g����IF�#�ۓѝ�R��+\t7>8 WM�vR��#��o���:菴���R
�9T�+�!½��-��{՜Q\�jߐ�R4��͈�Bex#kc^��m�<B����YE�uC���("n�K�~���W��z�̹3���z*��A�a'm�.C:��<�N�ݛT���t?� �`i�P��t&���������bȭ�D�[:���S� ���ҭ����[�N���}�����p�7���MZc�x����_ni�Jj��:UZ�R,9I�cQ��s�u�k&���sa��d�hi�N�����.w���F[b�'y��t�)� �Rr�m�7B�����JsbqGOȋ���n��<�����z����9��@�Vϔ�ʰ�ԗY�$Zy�����t��K�"�B�X�L*��H��}�7�{��f�כ����(P�)Ь7��8y�'�l��Vߝ���~W�}���kuhm�?��0U�'���ޏ+�cc�C�	~���S^��#>��ԋٳK�@��_���~����Y�6!�?ؗ�
ҽe%:5)2b��d���W&�-��x&w:�0#�5D9�E���.;���m~(�nu�1�g>�L�xg=b�Ɵ-���D����s)K�za�i�Du8DV�-���&���"avC@�U����5⣦XA�*� j�b�.t�����ee4W]�V���Y7R�?�|O��7M�n��b�
�p��?����ir%��B>���d�3�?K�[=��UP�;�c�1�*g���4��µc��F�E2h��%:�~"c�ލ�1�|a�7|��f�gs)���x�[���ܱ��F�|�>aC	�jՕ�@�v$S���g��d�z+�<���0���ÞNK��RgrXpF629�͟HB�$����q]ӈ6��D݂�ue�]j���xNw���z��� hT��р�h��W-��Eh�7T��Ҕ����f.���0�|a��y��E�/p����_��K���_S��P��&�_���uT���P���y���7�Ol ���>�"1��F�`;u���0� ��$�{�޿_����~�Ų��5T��7:Zq����l�u��¶sWq���T���];*�8J�"]��;h�o�0�����T,qu�&P�H������H��HC�տ�u���	��PY7r-����J��M�P��-8����ӡk�s.�D!��>�Fӟ	Mf[�! �f�T^QzE�G��.��û���>� �kt��ܮ>���(J�����_cRC��q��~:ry�a|&n�¢L��,�@z�����<�]���������g�}ø-�1boj��R�VTUi�"(����"6E�U��VP�W�Ԫ]�P[�M�_������\�y�{��s_�:��㋍	t���b�q	͛PMɇ�*���	�萍�]�jǕ�Ƴ��p%�@l/?�� ��D�'S�j:Ji;���}�?�>���Q�B�ɠ���o����U��[?B1���p4sL^�y	E��ë��a�V��i�^��,��C����}�Ê���H�k�"�*�JR۟������1I�#���H�#Lm���T��H�����;��$�fRW����w��;%�,ԑ�i��C�'��~���D��|��C�v���R�`_���r(}��;xЋ�F�!�
�bA�Ւ!�h�{R�4�1O����Gt����N)��p�̅s1C\w�|o�'��؍ui�o�������\m�
C�j�~<.=]��AF:���X�.�����N)5\Q��,��ǝ�f���]�&
t�u2|0Zψ��ԆY�;	��.|z���Țk �x�7��fi�Ƃ���ŭ�y����Ck��{9 *�mn('(g��8j)f��~�4�����l`���Pw�J�0�`�O$y�3�m��*#��ibt&�ʰx�]%O2��M����ћw���yb�")�ş�ޤd��U='(�x�5�f#���?}��Xt�A�W��n�b� z���[�[��P�����%��B�?4;�����%��Z~��!Z�*��� 	�7ݸ�%�%]Mg�OHH�� ?�ʜnL2@�H��tS��W����N\7`� &�V�/���m���t���Ӈ1��77h&Pb`{�yO�+^�0"����%�1��RhI��� b`� 2�C�
���W�Y����'��,ϳ	�<�L�4��C��))��!����7���M��o=5�o7E� O�s�M�ͳ�itVɀN��.	gסq
��RrY�P`F�wm�����=�O$��Q��E�g�1`F�׿�#��:����C��M9�Kl"��o���>�ƻJ?+���ɷփc�����SL���eE6k��Z'��Z[����v�'��$�Ǹ˔����S��8�u�S���Qps��J�Q�,S1b��!��ܡ�],Ie���Dr�&]7����2�V�S�6Α�r0�J2ӴFki��U/7�Vo�����U�g5�~1R�6�A�_�S�Sf2t�� d��^�7ގ&��o�{j��Or'��J�>�����>�^cC����ѥreJ���v/�2��h�V�W��7wXs�c~<�r�T��Mo� ��B;Й�iĚ�Y�yv^��W��8�@������������`c��Շ�����4����GK��d0��L�'$��]��t�,��K��9��a@�8Z��=9��kJ�2�3��#N�Iň��a�U��pD�ՐQ����G���������"}�EqI����	��vL�#��N�R��� ϣG����XK���ןɬ9�ʩ_@1O�J�{y���M�t�5���&�����70���3f�#�L��n0-N�4�e^E�Ծ�+�d)��^��2��� �Q�+�����F��?�a$�b.Z$�R�yO�x?~e�����h�bE��"���n|Z�E����m�\�i���ac�}c����C�� ڤ��,�	�Q8�>
��ȝ��B�ѣ��ؠ�r�?�!�L*x�/�fQ���a��p�$��+��r��i ۰36�jd�p��������6��.;7y���~���a<I����0�tvb�`���wDӮn�,i���iS9����:���2a��#؍K�մ�N�ѕ�ͼ�Ħ&����N��u����f>z�v=��3Ug�����$���p��?e-t��]�a�("�l^�*l�
����N͆�;��u����֣S��^U����ܧ��##J���@j͹- 6}(|�E΍0��1 З榫T,�b���L�:���]��|��H���>$�aYȶ""�;pLaͩ3��>eQ��3pmJ�q��ȼ<��O��E9��^$�p�>���ս��g�������
���
y#~s>y�M��n�]9��B�IVa>>��Q�u�;�>�oߏ"ǳ�8�=='ծ�\	�9'Q���9����Tֶʄ`A]�� p��n�|�p�&M	`�w#�m��u�>���uH�����ɻ��=F�h�lgS/Sp��� �������݃�LH��iV�IsȆ��� �*O���A	�}]ޯ�������=	�o�T�YE���2O���&�e!��;x��r�\@v�,#��{#pBx��~k�hst�R��UR&�1 ���A�J�^;j��O��;�tt��+2-<D�,�ͪ�k�1���յ��q��\B^�==�%��B\���0��j�fgk_\=��ט��T��:�3�V�K�����놟����b���3ޮ��s�Du�͏1����䴢)�*>�P����T�* z��4�G���cn�h30�v��$[��N�FԠ�{U�ƿ�Of�<�#��o�qj)�G|�ڢi�W�RWĞ'��3::�-�-�$�������k��U�d��W��-ŷ���$����-�$�*8����9̷�&V�z>���K8)�XGt�f��Eî�o��<P�C�5Ցfi��&�VSع0�U�2RT��_?����/������t�_�F(��Sx���s���+��'$d����E,��^��&xm�c 9'���.�d�U��<�n��w���S�v_~+��T29q�m�EK2'�PbB����QQ�Ȥ,q4��H;�w��4R��c*�\�9��G����-�o���b=�Ezw,\HG�fjf�=�|@0�?�%Ky������-��n@,�ۀv�"R�|Aq�ʆ=s��4�9�ܝB�hl9�|�0*1��	�&_��Jde���᤮���:tpN^��c&X�)��1�e��R�~8�n�G$�S�[�h)����VLM6Uӗo���+c����� ����gҫb��AD^ �T3+7-57ѫ�������llȞ�\v�����'��]�Z�N�mG�dx��#�_����v~��}q�$-`U����S��H�`
�M~�����~P����i8���#���٨��/�N+_Y�Y�~�]�(�/b��Q�W�٭*��6���������\Y`i�X�C�3����E���Cn��2�>��n_q�בS��ejن̪��;��
�G�ó����2�m��W�&u�KR���*�3�'����D��8���X����l�ώ́ߞ��m�����툺ߟy�s�}���zyuTUkfE@I�c�W�bW_���}�*q��)�&��ȅ)��nlM��=��N�_�|�u��E�?%���t�����s����BTS�V��	W;}am��'W?Mu��tܽ8$y�@)��;LV�}S�����w.���,Q���/��Wfµz�bt�w�����4Tʾt�-W훒i����x
������[�ȼ}s��%c�Ң�ƶ>W>��͠k�z�#a5_*�;�:���FT��Q�����*
���{\?m@�Z��eN�>��Hm`�
Wz���|�䶳��5�W4B
��1x^�g�Z)"�c�G/V�f#�
��Ë?j���|�ɘ�
��4
1�f1�`[Шr��?�������+���~��K��x�l���~� �x[��#�>M�;�o"��~��#g/nh��&�(
�#�2���I��HK�B���@T|�G�)������,��WQD�Z�΋7��X8c��l6��=�j��
��'���бJ���#k�;1��K���N*���E�e��EN�F"����B#�Đ`Y�	�H)���;F������t[z�v��_��P���H�+$�' �F)2a]����18;,��YW)p��3N�}c���$}���%���a�An2��(��\�>�a���0�����ᝨ�5�{��������p�
"+�{!���sƵ���f�/q_B�~���/�������E�$5�o=�R�U鳀�G		Cz(1uRz��^@&�U�>Hia�� �.�]���W/���_�F��P���wt��p��p.^筳,�$)�1�n�
����#��%�\ �\� ɲ��t��Zo^(�gUo����h�x�2u7�{��}̡��y{��o�%�E�F7���p}K��
��3.S���.�P�~*�!Άɋ1�U^��Z>��{q
g|ˎS�s>l��S���?��;��vA�ji5?g�#N�'O��ݏ�7�YR��J�K!N�H�҇]�k���\�4 ��-k���Yu=��Ծ����S�׭�_�b���	�2]y|	�#.�::���P�0D���G`���StxfG������O�_���w�[
ߧRRc�){�4+9�]urt"k	`C������![C�y+Q�u����ix/�7��z�u�ͬ�,�t���!:B=�s�}���y{�k�����#��r+?
��� ��KW���.Ku`w��/_yT��wުHX�E���! �񐯼���6 ��P���yј~#���H�[��G�e�u{.cw�<JϠ#/�㩖���jo@��]�!i�s�:�k*��px�E2ܭ��U�M��K�xV�?���;��y=E�~���9)y
E�v�ذ�����Ö�[���q-j�%k�NX:��u�����{���&t��*R�됳�N:-�9d�[5�V;��K3S݃��|e,��Ԁ��>�(\������0�O����we �(��j+$uz�5&W��[}���%���~��f{c��o~��3A&�	Z�����RNӉ�_^��]��<�F-t��:h�\���@{�ޜ�*��,K��4�Qd�U��qyl���o�0԰�^Tc=�N���:�4�K��m�\�\Zb4���� ��c�����L�Al�"}B`L�&^�I�>C�%�:M�K��#�Ȝ �/t��r`C��0�igZ��?��w][/������\�!,���Hn��&��<:��M�ɦ~��`�R�p�Ò�5�p	I�0Ӏ��R�&ӓ݇��,3S%v���xϚ��88iy#pL��Ѕ��� ���b��,����P��nѷ��&�U �O/�6��Ϥx��o�3v��Ǵ/ɟ�X\���I�9�j@k���T ���:���ugn����������<y�E@�N:��g<sa0ѯ�hQ}/��n�Ϋw�h��Io�N+�/��Y�ӕ"��~�m�`���¬���{TR7]�/��.!0U$�1�͸+C��5��(7����9�+Fy�>x�����@�d�j�~������`�g���[P*�:��?��;��~_kx ì�1�/�ٺ�����������eS(G���?�@��(�іx�"�>~�#�ށ)�я܄���Dv`��T� ��殁�2���;RIA��G�i�Jmi\f�T'�v�Q�m�2$��%֬�L�>�7�in	n��n���m�H��{B�N��a$�#����o�:�Y�a�/��w G��q:D����o��,*,�ʇC�f�?l�����R���"�͆���P
��>ۧ�"���c�h�A޽���M\�ײ�N����W����#{�;�y��6.'��Y$X��q���ٸ���8r0呰r�U%m2�䕭&!7��Gv���ާMS㷷/���,35���$T�~�୘2:�Op�T3�M�d&�����Ǣ���b�co4Q�L�,G��W�vO�My��1IvOH*G'Z,C:�כT��9�ByWA��k ����W,�΍�z����kx�ʄdx��W�Z�X���8i�v6��*��V��<�E�q����^�e*�X���)�>��#���2���-�ؚ���\��lin�ԧߞ�U���P9���`R��(#c����/m� �9���\��6�p߸Ԟ�g��"�yt#dO����W���u̩��y%Z���_ݭ;cHJޟ��fc0�X(��7/9���X�~�͟�RžU=�+^yg�*[.SX�� O*nv��w�u1�a�`@�k�z��~�z8��u`Rs�I��}NJ&g�8Ǌ4:l�Tfi��1�e�%��6��N�R�.*�5�OO ES�1�� g�2�eS�9�M�z��`E��S)G�|��]��}}W<ež�Y�~C�$��[�JzA�g�bGS��ݺ��cF�%�x���#
nw-���a���)�	��	e���n7Zv�&�觉@%���^�xxGɋ.����F������Ȍ�	�EA�5 +6���5�<O6d�����];�3wCHJk�W�?="9s$�e���Ħ_)�~YNq\�> �����`��Ecc~G��v��5��2i��v0��� ש������,s������Z*Z&�ᱻW�4/�<�Q�bVjr�ͭ툹ܷH���AJj����Dp캀�,Qrg�}	����m�Y�	:=��5Ԭ7Pb�'QZ�^�ʣ��wb{p�z7Cz����0ob�x�)���r�}�����/Ee�h�d�Ov��6�ӽv�#̀<��|I��6Ks�Q 1T8�#�wG+9�8d+(i�����l�w�����sS�pf��KM�3d�yJ�cc�ӤcI�7�ǳd�W�x�0��<n��g� ˒7��'�� �'C�,��jVg���� P�U*���Wu��b�>@�3;�N��8���_�t%�Q�̶���ɪNӑU9�z4��Y�7ZF��f�x�w�*���}��$N��Җ��� �+3~�7��#$�!��2B:��W��G/�$��wŔ�� y�3�������G������[=��e�j�Rg5��|�!8zv?n�4�fz�1��F�s��s�+Q��U�G���0o'�����	B��!��t���ۨ�M���6i��6�0�����@�J���`_^/1>��������yx��Uv�2�i��FI��z{�v=���6EG�$X~�ߗJº��b_���l�����<��+��iL8���`J�Y��{a@�M/}�S�{I�\�ѿ[�},b�ʔP���5:0..��Y��V��%#��S��u��zI�O/�������vU�SD���y�~&�����dH =݉u}f1�(Q����hއL��҄Ë***Й��+�e�u���_����舊+����O��g,1�����k7�#�2K��7�+�}��A��T�J���5�m�*!�"7m�g�N��B�p�E"�Q�w2��ݫG+oR?�OW\o��.�ku<,�[�j��J��+���=�J�&n��Y�7��p�ܝ���oZ]�;��qU��}_=��~[����Z��P�Մc�J�Z�4���t@b���h��%srW��|���>G�k��L���6���BIa?��Dx�fc����^����l��ڶ4{R(��\��K��wv�R.CڍBg%n�.	�B��Xm� ����Y��R��W��;��H�'j�t�~Vi(��΁�'3�DԘ�5�n�?Y����ȃ�����Q���i��Z���c=�s���O����;�H4������%������ϧ�<X�x��z�d&�H[:6�q`�u�(�x��RC)U���g�J蛧�@�:�ϛÁ��v��z�V�?���dV��|⎫\�>�����s�6� ���C��0��bX�{@bbl���a�HwpB��t*|�ǧY�䎢�C��_��mr���-���.H~�� X���,MQ%�6`�������_�uOj����vl��Ufa�roV�P���z�2a��eü/x���|E�X�kץx_;ᐧ�7W�ְ�q��)Eg�s�ׯ0|�"�W�[�7�U|��˧����b�]Ֆ�B�V�i��&��AiF�p�ً3�, ���(S�P%�)+28���2�`��{�N�	��~��d#������I�$��>��heõ,\��R~�|��|��M����f}�^є��lQ��Я����b {��{�ܙ���S�����O-eߎ`&z_ewe�j�3�o6�d}��ye��?;�����m�+�~�$;_��͗F0/������a����&R^�,e=m&�E��Ye��G��c���S����՟�{q�`Vș܁��>�w��'w�5���-�F�I�����P�=ԛ�=���l�R�wr��!�I�&�y�?R^�1ry�Y��P=׉���b���s���� �f�|���^�e��/�Q^%5W#UB/�Ҁ��i�T]�A,���Q�b=��[����#�O-��Hk�e�+�lX`��6L�9`�;ޅ��0S?)"i��l�X�9�XI�#y��Y݆u7��lӲ�t��@�(3'lu���9�Dd1`G�}F�~��OBt�fy�w�H	0��,r��i	`�$kPp�Y'�h����C^⏺U����$]j�	/�����k�wų�=����3L�=%��7�����he,dݗ��Ч�%�a��r��ކ���e�����؏��HVx4W(���V;~P�qbϴf�Fe���vco�se�Q��-	��C�F>�ƶ�Oe���X��X��ׅ�3�)rlg��N_%�Ao��8v���777;���]�s\O��k�><-+���	FR�<bE���,��=����爏f|ʟ ^s�?Cρ���B��0��6��M�fM`�ʱ�#� ��˦��m�Z��2Q�-)��S���]�W�ݗ�M%<Oc����nf�l��NR��	����S �1����ZA|.�l\cZ��v�O��N����=x]��9�/���vqaJJ�eA8y&(�-���x ���t��������Q����_s9��J�\�|��n�R 5�ҩ�Y�F�0�aQɕ����ߎ6���@�Uz02yujF����{�ιƓ�7�w����y����VM3��H���Lp���sS��'CD0��wV��wk���'�\Ujb��0����ӁH%���2���R�}V$n,�FO��.q�F$ƾj�ч��ҭ�������-p|��/�2����X�D6�9΁�)m��05�|߄0}ٮ��	�� Z
Ĥ����Wߊ;z���>�xѢ�e�5:j}�[�t�V8��+�)ދo��E�C&�$p؅�Ǡ�:��������*��-PhV��K�HA�_���te�_i<��>/��h�L�ۡ���\�� H�)QH7�O�|l���n�����' ��nss�_w����w����+v��ݿ�P��OA�v�q�2@�l�{R�����A�5`5��5��P[��.�tm�u0��e�iUȊ��Bm`gO?��jv�"�s?go�[Z��֮'��(pNZ̼����yt�y���!��"��Cf�>1���]2nx�?�y��<o�|q�U�7��X魠���*�ri��D�=.�9W�vpz�q����搾S�����T��_�F�����l�.�����m��kR��b	�G�~2�a��|��]�����o�b_�_e�t�:�����V̼^lȥ)���V,]������ŕ���A��/C��מ߯p�QJ�����#"N���[�;*��H�JUl"X\}&P����D�sO��S5v�qtu���l���SN�;�ѕ�D��}�m���C���)Uu���d_��&�LK�����4MhK���d���㫡��x��g����sY�o��,*׳�wf�m�bQ��a5v��'R�i��=9�յh��!�d���/��!?K�}w<p軻�q��q�82}����~7i^4�`��h[����+6��
�j/L�����",!9�5r�u��m��w���<��XU���z8K����F4>U��f����-,"Oc�jH�#�w�U��eapG$:��ò=��^�p��
�RSI%����b�|v}bA;��a�-B��dP��X�R�j�j�eq�f
�<��Ǚ\�S�� :ŚR,rI�:k��X��Q�j�(F�Y�˺�u[\t�p�-���U����	}6�٬��ǌ�w�=K/��������ŉ�u��bb��"6o�	s�jV����!*Z��|�ZCē��虱�������i�%��r�J	�k�K���Ŏ�oXN��8fw�������i���9�{��p����on�.$��x!S#Z��Á �S��-�ÄNf�)"
��]� i}3O�W����B���3��e ��Hr5�~T��u�Md�R/*�	Eťɥy�ʥAS����{�9���k�M��W��?'����tA�~u�0?>��#s-<��u�g@I;N���)u��^�0���6����uHB	�g�N�)D+�s��ֳ$�5��rȢ���h�{3�T���4�]�0$��D���T͍��������J%��=7��h��Z�:^8J������B]�
vXb^��K(Ѫ��{���� ��t15�U�)�9�h
7��B���p�[,�#Q�1�0y����r�m]�{k��+EjM�Z��-Yƺ`Dp	��xC������Ak~�i}r��Q/���2��&3�d"�n�z;c�.����~sH�yq(�cӋ#�:6)��P�N"jk8�M7� ��QN�y���S���9|�d�3�3!o�Ȟ�@�ܾ"G[}TDF�m�w��/�G�Y��"��6Mm�0��I�I��aw��=�;9������F���Y�MD@�3�>Ȝ�FY��҃dL�g@s�c���h���	�7m:��w=E��_�vͣ	�+.tj���#�*�W��1��u�u�����#/o���� SF�W��h��6/$�=;��!\�:��^}���7�ҷ�l��\�����O��*�&}X���	\��S�s���t��\�y��؞�i`]�[����8#��t�,��N�K��an��y�`�QSDK��|p�_�7=�:���'���<�I�9��7����6+�X~^��`���W���h��C04)IU�ȃ~E�	Ir�dP���!�d��gpX�S��;�b��"L�#���,�so����B��=� �pq�gS����O��P%m���?2R��A"-��w�Cv=�?�m�M�EG%2JX��9.|ԩ��tw�I*�1���gǸV�즤<K�l~���w�q������l����#w��/��,Z�s�\{O9�<7�,�<قG��+/�?3׆'e�e(&�N�{_�[�kOp�/���p(ů�}���(��֍�G�`��n��]����lWO�(�*s����RS��%xcU�ҋr���zWʘKҒ��������ރ��D�m2����-�if���4�y����wx�I��ޥ����(�Z���7�y�{>�n����u�-���K�4��=�[���5��{|k%�<ެ���V�����a�����,�}����=��kiTܑ��6�<<a�7��l�����N�?�������nh^MĒ���G�=�i�Y��mv���a��LcQ�O�Y%)���!`ȣt�U��2�Ɠ��<��W!�<���C�͗a<y�^��ɷ���p�QӇ5ّ�Ȳ
$�_����It(�~�)�%%n	�Ǉ;�ʣ���E)��$���5���{4�2��b{M|�v�lk"Ī�,s�Z�1��W��b�cp4���'�H���n�RZ%�c���1Qƨ���,e����8��K��N^�˕�;h��XI�ν�K�'1�_�R������M�w�#u�
�5'��Z�y�]��!	���ɛ�������Q��(���Ki��W�^�5TLm��d�Yqn�os��PBLq!<e����P?�hQ>�6����~�0>��@)V�����>�Av��K�+���&��3�� N%��^V��)�R'�mB��܉n7��P�(Ε5Oܷq���?Z/�g�ݍ�R!�\S�bQ~�1�]�X�}��+�xvQ���Ţ?!��kKp��W{����x����D����y@韫��Z�B�?Q��k�����Vo
o4�U{�z��\�a�7�䯜��g�	>j���2���(�wٗm�I����gEW�;����E��p����6-IK�x��u�R�Hɻաu�%�}V� Y��7J_CS�`L���4�b��jjyΛ����a�oֹ���p�y�=W$�m`�_��+�r�3�g�Fm{ߥǜ\۬g�t�~灺pP�`�qy�z�x����bA~J�k�����G�/ZONc!D����٩LM!٬�:��9���&��~4�C�g����匍�\���[)�M�%����	/���h%�ᄣ��"�ž$\Kl6ό!�
ƞ�:���awd����4J	�r�7��u�;���T?��3o�o��[u8}|�A;ѡs�aj��p����?�t�� U7~-&-�ow�W�$,��3���>�-C��f>�}�3֧d`������������6��O�=x���b���FYF��.| K�s3uO%�v����ݙ�x��Ǒ�;w55��@������+�uF��FAeN��;5��4f.� KV�s�<i�C����9̯�����5G*-�tׅ�Xu%�d�z��#��ޔ����$�>��|�´咿zW�k������	ko�'
�WkɛAW��|���5��N���+�_��پ��L�r�Ж�6��t5[P�adq��Q��t���q'�����e�U���x��ڎ�mXԊU�D�R�������K�U�h��(�/H�I�o���n(����%��hd)�ă���g�hc���Xb�U��k�bfjd뽿�T�!gcW����+��ؙiA�t�ǯ ��%��˧#�?�Iŉ�E��C��0-�g��]�_~��?X�g��ंoQAT�l�S+��\����Иr��R��������g��� ۦ5^��-Q75Λn*ѧ�i��w���T^gL�B��|fq�����Y��2�F�z���|��?r\z�}d�[��0%��lOW6X��3�y���ґ�
�}w��H��e7HtPP�3#7��h� S��`��=��G:	��#�i����@�����<y���;�W���sV�0An���騰!��[k�L�2!�vR`�1�Hс��~��J��3��\�3���Ep����l����mH�T��O_1��ʵ���zf�\R�qSߟRX!y�p�̕NP[��%��%���$Uޝ u�iX֟Z��@ ��K �ph� cQ����H�c����;U�c��y�u��L�Gb�k�1zddҕ��\%���qsVIeH��DQ�*>T�旑a�+P�Ý���b�#[b<-�V^B�
!_��Q+; ���&��b!K��X����i7W�R\=!4�O������MÈ���<-��?��� ���뭂_��ȆOha+aȜK?�3A'�-}����5ᜑ}����]F���'�aS}Q�Zs���ͣ��7��������b��f��F.4Q��kMj���r�]ǜ��$���"��n��e@��j�t{j�4[?��w��·��U�]/��YNUW�кg-����g�\��D'�be�������E���$A��t��HH�98��
:��=ΧKy��:�[(K׻��L���W���r�(��ͫ�!;��猨?���'� �%�tD�C�	��/.��������}����RՍ*z�"�%��7����Jx�'���'[����������<�n:�N�������I0|6��8�K�����H�qߣ,tY�];���#df���ri�^�3ފ�sz�c��פG������XYTl]����MU	��x	�sm�����e�5ۭ��7ޅ��P��дa��@yy���i7-MKy�|4n{ԫ�YdEF��V���%mH�/����ߘY�ˉ�
9�,l��h�C_�M�k{�pKXs3-�c&�D?`���G���OD&H�7����V� h�6u'���Y����z|����Uv��av��`�,�.���ٟ�eA�
6������y�	���eՅ4L�t �C��/5$i�oB�p��,��4? 2�6I'J�ig9f�p ������#�*{�|��~�'�&A��i,�i��S�/�Q�s����0�(:���@��Io��Oq��;���u\����D�LØ�2*�����:�s�+�$�3(�X9�k�eb5��c��ߟ�Z���MՅ�!f��ϾeW	����aoE����`�ڌV/;��'��]����� >�ZK����d��͜�BTqB�;4V=s���gYQ�򖁳a��Nk7�-�=�[zz�������N��~^}#�DıOl�Dar�N�b~�6FO�T�9UTZ����2R�h�"�I�d��5�l�1�x��-g��q�t˗Q�H_����y�ի�8�#P����h�GsTW����� k˸��$��su֜DK���s�����T
kkwv��̍z3�s��J�P�1c/z��GR�㿼AF�%M'��!�fa�4��pu1���]�{��'8�OըnT����_�+T05��v�c�|�M�_�f�Z�X0�ԓa�C��a�QUgA�>)k٪(F-�B�������������A�G�����Bh!�8����zA`,<���Np�Ռm�L3�I�R'��2:�<���%����9Dۃ�F��e�Q��F�{��G�0�_�����=���`���&��gսs[F,H6֜��I���(ң۷��m�����eg�i��ÿ�*ou�XF��lqPz�zd�!4��ZGx�� l��K^sqki`%�}�#�����@���p��'��&��}�[�*��
C&�0�f"��4�Q!�L .�>X
��?A{x"��2�`�w=4P��I���|}��yJ�'A.�E.%��9�o�"����QTϊ��2$���7��U���|fO�:zl�$��B�xo�������_�H�OW9��,�x���&[K[+�œ��T�0�c����Y��>��� 6�sk�o.
9E�r�y��Q�F�lfb�@/�]�=3D�&1BR'������p0.�	uB+�,�:��17l����jO��{;ﱷl��"YCH�n�WI�}������ޚ�]v��%u�6���q�`3�8��(�Ih5sμ �W�3�n�#����>Uc��0_�!n��v�~B��P�>E�A&�/��*R.�}��@ie���F��6?�4��Fr�<j��ٯ(g�Em3��`�~3����QE��H��i��6ap���ilp+-1q0M�tC�����,%_���ڏ�xбn���
�|S%�	������y<3�|�'�G�vѦ�u ���oD��z��b��%
�!kVl��Vp_X��l�_�n����������58�UQ~z�+!O$?�TqG�'�i���4M���/#���BJ�Z1K��e����$e�Ї�U�Q{N�v�w�1���c
H/��zZE�3�K�Й�N�g���z@:� R��4: >��	�&�*�����-|�;5�j�C�����r����3���p�i���X_~KzϺSk�H���,�%/R�o,2��y�?d��&"E�Jg���D:��o�b�V�&Z�1�J���=B��ڮ���k1�h�,���U��N�$��8�*n6��d��ȋ��g�b"�e:���t(:�����Gڏ������:��?3�1�f�\�(:D-e�]}���/�~�\K�d�얂G'Yj�7��0���jϖ��2���Wg���zg�N~W���Y��wnrJ)����(�q�*A�J�^�6��b�P�9�S$��2l6��,��䆛�F�>�r]�]h[�.��zE���^����;���%�`e<���P�Y0;��0��h5O+ˇ��{�:I�9e�"q�3�)r�8��c�e� ��`ҀV����'1p�p8y8�;�54G',$a�!�{�R!7}y����
c��9ց>-d��[+�l�J�	9�^ҹהMb��B�E8�����oЫF�" � �Vxk�b~#r�&W_���4D)w%�,_�%���/�ۯ*�@���5�Y�y���|{����@�&9�}l�)#��[+H��6���E=�]@���t&���ī6;��,����n<PO��:g��"֋�;��
��� ��x�ə����f[o��W�U��K�&�����31w��/<L����Pf̸4 W+]�.f��YdVh8�d���|�V�mS�ٽ~�oDck�@WR+:��w5���yƳ��mܞA��{��޻�*Q3��75kF�nKQ�j�({�B��]5�"�h�������<8�s]��y�������I�\`�8^�X*af^ai�	z��� �ܢ�/AI�'�YX?Or�5�����O��*l�������n�|��K�˺˒E�<������x�AK��;=@�"�ZWv���}|��{�E�W�ŒHlI�6g���u��U�7�.�'�X�!�>�a{-�(Ĳ��;���9���ι���э-��*�\���e<*�0f��~� ����������͕�oU������1'�:����R���E�3-�3��|e��QV������T���Z�t=�4����&�J��l�F�D��cI�� >Tڮ��b>(�?d[^��%�xK@�uJy����B �I�Ѧ��d�C߻�.�G,��@��Zm�d���0�����ʋ���nSx�r�� 9A��Q0v�U�[�.Ϲ��OO���)�ݕ�ayϙ��gS=��N�K��'�̺J��#Ο,�g�p�\��ac�YS���$A��Ax��4⁻�v��3��t67�����c8n�bt.ʧ@n�d%疰vw���L��%����tk��r^)��'c�~����e>N�  Ǵ�N�KtW��jT=	��|��h螸�¾��+"�n�3�q*���y�A�k���ůXf��Zk��(+�&VM/�bU������ȋ;5І޼ `��+��C��� �d�:'�����3{r������#Zn��(�O+��{�4��q��.4G�k;.e��4�r�C�0xS䋫|�3��Y��|�C������^���w/m�N�%k�׬����Z���)~��V��r0�����0i|�t ��m�~�MЦ��O-sF�;�J����%� ��A��퍪n�V"Q����sR�Cie�٥�)6��d5�Pɮ��y���r6�x��*T�+��	7y9I��7�q�3z͆�S\Z�O�'$3>}�P03D���>}IN��V���H�hmQ������7d3����9%��{������SG���~yah�H�
PSRB�"/��j��WIU�TL�M�D(Vd���]Ա����(
o;���$���mHM�oN�G���<�I�8~��AsQ�2�{�ݳq�]@������g,�4`���I>H�$\� Vi4��}����t��Ph���Űa���1!��X� �C�����k��H_r��������?�h��M�]+���}�(r��ROV���?�TX�7Ҁ�V���d�������������W�S��!��ٳ�JP��	QZSB��㬄DgAN�PJSPz�9�v��9 ��;-O�R<A,�Rn��T<1�Pq�R��W�u=M=���3
>�����ep��!bɬ]��Hz*����	Œ�By]v�S�	��Y��lNv*W;/q�1���urh�Qȼo�6����yP��ؒ20��L�DA�>�.5W5�^��J��9�TGɖ�u�D��4�i�3�ß2�6*���>90�t��9������CJ1/����������|����>&&�k
8R�*%����]�����޻Μ��Xd�=�X|��\�\\����J|�ꘪ�҆��G̖�2^!���;Ac7�:�"�|�,��_�����E��)�g�n��g���h�65����P�	�ы9W�)������ �� ��=�>Z�C{�6�QZ,��������Y�C�_oT�6�L�s���,7J����f��y$�E`��_[�GP<G��i��_��L�f��h$Yq@�8͟���(�aƢ14!����e S~��c�Ms:��3��m�2#�?�z�ӓLMs����W��R�j[H؟ ��OG[�i�̀��8bMo7�R�X�e U��b��sVg����h�:)���.;@��TR��J��������1��d�Uᣛ.>�^���"ä�Q����I�D������xL�M[����R"q2]i����0�BRo��<(�=b�$2E��#���PdT�{^F��j5,��/ 3N쩯���ށL�>��ؙ��*�T�v��?���}��d[�vE0�p�CG3�姷���M�Tn�oez�(�o������UVt'N��뻮�wwUx!� �. ���-���d�����)�j(��m���{�U�tT�q%��oS��?^�/K��kNPP�!��%��ݿ��o��F޿K�re$�궞E<�*��&�iKH���CUE4�ܥӉ��9a��	V��"���Ʃ6�z�i�ϕ�)$�0�<��?08�O3��<�d����K�6�oG`�$P@Z^�3<#w�s�Bx2yϷ�������l����J��t�Q�s�<P����h�>�J\
lexI�^^���uO���0�Ľ|\�Z�c@�>�7W{,��ݍQ>i����މ�Y��V ڐ�Ջ(�O������-H���OG��lsr�I�2b��#oLsr�z���6����񫩑����ƚe ���ԈOq���s���9��o�s�L�D������k��3��<;<�9�����qύ��-��AT�s�j��c&M"~$��a ��K$��xI����`V��@r̿���1`{p�2o�pz�W�[Nl�%��@�@��K@�8�k�KY�#�i �p��]l\(��$�/�%|��4�U���&���p����:������:Ϯ��B��"�&�w�����d�8����r�&%)9���s"|����NC!�4�e�;���\�[��c�P@���д�L�10{�ף�O�e�O�	��|�H�ш�PV�%��;XJ��� �.ǐ�8 ƀay�I'�'��,�&/T��C����Bk_�L�#<��ú�5H�� ^�f���Ƿ������wD~��A�0��К���kM�'9n?/y �։rL$�Ŏ�;�#�շ��.x\\`%J�O�Zfa�N�e<�ݽ[yc�H`���k��4/�}��#��A�[x�ۥ��t�䕼^�L��_���$x���yme3/�˳�,\'��	Xw�e�tJ��"H����ّ̅���9���)i=r��`�(*@w�p��W�uu7�XdG�3��s��kO����(�xN�h��
랑���ss( �P����2:�G��E����~R$�D�L<���MRa\���M�����If]���>�U�H5���P޻@�,ѳ�L��qs���	 ۯ5p*v;�c|הHl�����L��#��% K�X�D��et�� ��#�E��VI�>��a0�Q*�����1���@D�5�V���������ޚ� S?���ӄ�deG������$�"__x�G��o�&L���|/`�8N�өy[����w}�a��v�XTD�LϨ*�j����@����)n3��p{��<Jq�ɧ�pm���K��������M�i���E��#W����o/�*+ص���D<Ѱ����ǕGlnF�p���JI����XY	|r�,Ɯ�;^h��m�1l[z�Y�E�U��O%z<����s���$�JE]m����w$z�Ve��)����H����ڈ�Xk���u8͐�Ԯ��u��o?��f#����*�������U:p1zi�]z��G�J���"�"�,Q�����{������jZF��$��)p`OT!�?����Uֵ\�s��Ny�����t�Ԟ��&g�ie�g�J��T^���sfY#�8귮$�u+�{�~"d�%����!�,(���U�����(�8u-����Z�u��i���?���[���E�2B�9k\�^��	H�|�{�;��
���.n��~\��?�2����[�7��.or�Mm=]��D���_π��,v��η����f,�(>��yW��ab���t7 ��)�q�/�￤%m�ۿ~�`W���c�?���0����t�����1�W��D�r�����C�"R��h�m3!��>�3�u��
V2N8�2�ĖR�Oa^JG�
O�����7r~�����J�Apo�IJ�eP�X�����Ӫ�4M=2v�u��E&B��8��p�����,�RhH�#s-�H�F�=4��sm�~�͇���ݟ����|<fP�}o��y0��B��v:g ��Ӗ�<�]��蟹��sm��Н�fʳ-���4~�HA���W���@��K�����5�q��|��W-�+'!���ib�e�(�Qd�Ƌ�3�F�{H�E�hP�y̤w�������a���D}�G��WѸ�r*���K:W��������)���5�9��Ԁ�����+^T��Ά�zЗJ.n���lȵ{�<��XF��Frh�=��\q�vD�Z�2�?Ҩ�aM*Bv\)D{�U����6^�3_�i����9�7}_��G�4��5���?r	��2cK���{�!o���>�%EF�#���6SQ���}+�}JN���]ͫ?'mi�J������~���@E���͜7f��_%#���u~��W�kSW�2��- � \�tx�9����\}%��F����ۯ����@���ş��*�՘'��4 ��ͪ����w.�f��`( ��f��e�K�K�(�zK�x��˹;{�8�ik��; ��� n���&S���[vӲ����ƒa_��g���>�7o�I$<�z#grYK؊|�2��aH�CC���N�ף�� 7�)��� &*�l� ��>E�'��s���ШZ�{ph�wd,�$3����+�v}B�/"r~y��$��]���%�B�g~hD�ۀ�H��-l{�Y䊻cR�v?~���Ϧd������JߔM����\a�3��� � �х��e�#�ΕY��i�a�����W���wvh r/��C{�Y�% ��Ԝ(~_|_�"����°Fd��֮�J�I�2S4Y�H9���5�k|BC�[�:�M��>s/��yAnV'ݼ��R���t�u}\�{�o�Jw����an�����DA�^ź��T�}�����AI-�Yh7Qeۆ֔�X�a���Ͳ�&rMK*]0�;J&��	���(N�g \�zMa�55��pAaV���}���#ص2T�­8�{Bh�\q����أCW{F�[/����X\�;a��X
8�$�S��
�e���D��"eGR	�X�����tP��؞�k���ʴ�֒���vs�{cܴ�H@w=���~�{�����j�:4��M��%���?�����?�f�˼�pikrx@�&}`
�-�s�+�xESa�H��H�o�f�ۋ��D�+]E,�i��L����'��h��~��+����y�M�, �qL���Qz��[���tYs%��]�D���g���g��ǔ�{Pמh��[ux���&��^��^c�J�(D%ۗL\��jD��P�;>�{Û����W�&����#�Px�ڕ�U�ZE��7�(x+A��%���O�M�t�?��>����ŭ}}�/:��ՓZ|�nI�����]'�h�K�n؊2���u�KZ{��;>`e��`��>��N�`�ћ�'Ҁ�u�����`� ,	���Ղ��2���K�8u�v����m�\��?-E��l��?�P+Dn3�}F1���|�`��ݧ� �>b���MTV������_�E*a�Թu���;�i��݁׽����R����+l����yX�*��� �x��G
F��̽Ч����=j)��J"i�h��}^� ��o�朡�ƚA}88�_|����{HÙ% *���V����Z�E�@ܝ% ���u�aH�@���aPoZD:��8.�d�Hx�XZ�SO���=Բ��]'Sy�]L�L��,��~t�}�֚�zw�Ze/V&s}z\����F���q[��� rN�%Fq,����N���qb-;��Ư>҃r5�=��$�O��Z�F����S4�R�6l�ci�仹��#����n�K���Ka��K�L���|`�'�̈́�[B-%Mo[;I�:��p�L�M�!�M��g�|^ȥ�$�k���xyt%����rL��w�n����#���� Ͷ��ۋ����s)S}jɥ8�E���*����ϥ�9����2g�|�ID4G~��R�ř �c�I�<�A����K8�p�i3���6g=e���������~��T�%i.��.��dH�B�7���Cc���ܠÂ�A��������
��5 �-,9�G��#n5�2��#"��]{�����a����|��H�8����ILNV^��X���=����f�0(���OJ���"���a�������:��^�����i�OHchrE
��ᮈ����
"����KR/������<�Ht��oVf��"�|E%頁��
<�35:.��~����g����2����9�,G��K��U}��6���%�}������-���{��E�`dw,DL��`����5`�)c������^�����$�?Hr�e��ov�?_���#� �����H��V�%����+�t�Jp
�u��m�W��i�Myr��Y?��&��Hb�����8)\	��KX.��,�$y����B��6Ad�E?cü;�S%ɀ]�7����J+p�� 5�;x�#?i��Ł�/ƏF��WȒ���p���e;� ��	�n�P�.qz�%~b4�N�1���
z��i�I��ѕ��SJ@�0NDg��S�u)�䗞2���2��������O�a�Q��Y�,,�Q'�I���Q,�&B�@F���{�Z4���Λ���aVdl����l����Fo�c���*,u�������&�H�+o����Dx߃7==���p��<U��SO-X�Q�꤭�˶�T$�w���7*��9H�����<*��C�n�g �#���/��S�9ߏ�Y��������������	9����2:���'��Yv�C�Z���sm���=�����"8��Ur;�v��������5�.7�<�v�_5��m�p�ѳ�2 ���cS��OP�^nl"��R:��g	�w�P4}$�4V���u ���~r�_}"h�M�o�`��@,_�{����si;
dU"E*�A*Z��&��@y�|r�\7�m�Wg/��?�_^�:ǒ��e��	��s�߲����	89|��AM���\�h�3��˩;"��quj�,�������Ӣ�C�t	_����3���Jc�kN;� z^�4g�l��
�"����6dz��9{�[�2��&%�7��&�j�S|Y\�p4&5s`|C�!��դ8y����,���rq��՜ss�����J������b��D��l�J�yZ��%�a��,�z�/#w-T�oIר�"�9H�a�b$��zn��6�����H�_��<]����Z�K�'-�\ZfK��uj���(]����ϛn���[���+�tEg�MB,�°%�6�sC� ]
�g�\:{R�-*Y�_��(l���j�e��;ak����i[;'opV�*�a%uM���3�&0��+�|�ڿ�>��������X�O��`�f_ϥ)+����������G���i8V����)dQ���k�]+S��z�R|y���m���CumL���wgT�sM��&�:ܝ���7������~~�P2x���0O� _$m��G3D�Ę���kZ���	s6y2�kFk<�رm���M��2�Y.9/��Z?k%�:G�c�HH�]U`B���և����C��1����w���z&�T%
�B�-�5����Hxׅ�Ʌ4����(�0>M��EN�TWl�xW��iR�=?g��� R"(�g͊���^�t�$�J6�m�:���=��N���K�?��d�$,S���BRg����N��hA ��HN��@&'���D�ɚ�~�����V7����c�"���O��hz�Ss�!Rnq�k�p��P���S)����3ђ���^*Mz<�%Q��hh�	��#�N����al*�w���ތ 4.n&�Zw
 �D� �ɩ��{�P?��sf��i3���ta�l���q���q�FWw��ѓu���fgۏ��]����� /�s�XN�N���D�C���+�^b|��5�%���1�5�Ј� �D%�R#6GK���#T�cȻ�<H���V�AU�I�/�{��*b�]7V�G��f�ys�fH�l�^P���V��h:�%[��E ���0�>I�7�6q��y1�I�Q!�Y^x��g�I��s�i�s�'Vq��S��񁐃�ըDH�rl����d tI0A�ąu��s�ZX;�7�)Ky��i�����u����~��fF�}�oR��i�Р<nYן�oѴ�q-?��j�2���f埘��r�K>��d�$��햞]�����=�V�,<{��;���?��mF^�y>W�3l_�����_�TV���T
���0���H�����߳
�
��~o���m�|X���&���l��Un��칞���h��:u�<�a�R��\c��y.by]ߘ��>�2����ӻ-�Bc�x�s���
K�;U���;k���zx��gNn���d����4s�bw�\����?��ͽ��������]Ë�;���}z)~�A|� [����Azv@,Ky,^#�[`O撃A?� ��`!H�M���9�-� �st�Jq2�� .���w�It��.�H�1���L
<�eY���=�<�/�}�Y�]0�{S�Z�{�^����u�n�iU/�F`��n@K�+qGK�`K����KA1ƀ0�|`.L�](�r�xu���thJcVr�Zw��{f
�F�b	E���ڭDwVH�3����'ÿ���"G�bSY��W��X�G�"�����v:Ϟ;�(����X&�"��ʅ>/8!�nՃ��7�T����f��� i[�r���Aᗩ�<���ǌ��\4���>�gYJ}�|��&��p��,C��6�G� �f`a���n�j	�tɃ$�X�������mK�}�K���l7흶I����\�[�i]ٔ�gM	c�9��D�@��[��ΦVM��I�4�C�I.|	%m��:G��,��r1�pV~w*����T ��/��c8HИ��Af3*gc��)���GǷ>���%L+D����u�EOlp�����T�^V�[�(�uJ���d���i����ñ�~߉��WY�G�/�[K�:_g�0��	Q�>S����H9���6���>S�p�O���I7��|.����~o���o��O�Uk�����č�]��+�G���T�����޽�jg��u:�n�����Z�nmT7ܛ���f��SK_;#����s��L�7��O�� ��:b�*\IQS���ʓ�`���&��Q�ЇQ��NW���?V:X_����Tr���`|x����0ڕ,P�d�l���7����K������:�	Rb3u���+���|��]b�-$w̓�w)��á�>V�e"�Ɋ��b;��d^|�߅ON�E���6<��>�&IBhٙЬ��4[�+"����_c��Q�E���#_�'KJ!~�LL�)x�������nEL��*�h�T�<����l?�n�!5畈Z�<EK�)��xt<B��YqI�U+F^��������!޷!�4B�kj�J������Z؜�e�{_S�Gp&��_�x���β��� r�^�d�%Y�Fy���J.Y��=޹3a&��2'�ome�W��v���B��sIZ}II����*\�k<�*�y �Δ K���d.�V�eN���ɢ8-!l�c��%�!���_%ӷ2D0��iae���,�Q'�N:�������7Q�.g�İ� ��O����Zo�D�GeO���j�
?(����(Xs�	�/�ʧK���,h����z�A�������D0�}�����B���5������		.F�����:�^4-�KT��f ����)f(�d�d��@ħd���0���}����;��1�$�1� _V���*�)b�∕�%)�!����S@�+o��1̭�m����'U����ǟ��-j����3����:��[ ��Pi��������4�������l��gY��
]��W���hDNE�wh/	d�}X�\%n��f���n�j�ne|'6����|�K�����s�ߴ�W�^��}��f�5ee�r2��kӫ}0B���D��K
��%�Q�n<��o�J/��K�{��c�2gd~3�J�Y�7R�-�����E�����鑄�jSb�E�=f_#�_I�{��g�����( �jߢ�Jqwx����7�\���;FD����w���G�v�`(�:��c��nb�6��X�=d_�0�u<Cʮ-�6$�y�xwt�eӀ���0h�Ǉ���(���f�����z��D]갿�T�K����a4���A�O�Z_W<y��=G���5��[�[��IH���=c�`���ZR�L�����'46���O��5N�,F�`w���B��W9S�2��'cv(�F�҆j���'-���_5ZX:%�gΆTU/��S�ǿ��I�Y��	�'�`�}�kzEz�� ��sca���eAn���BGH�<n%п̊'<+���f�k�����I�1H��l��0��<qfJ��r6)����g �������:����L��:��Rg�������P[�����-�j�U�&�[���"�f �� b��1��P�/�ԕ�C�C_i�����O<��,I%�(6y�wɅnf�k{;�_�=tJ3ݐ�1�N��x�m@���[3
�	�{G�_��7ԽSV�N\J,��[�[i.�\�&iĠ=�x�B�(��N_����Z��"g���qE"�����T*l�� ��^:@��F��={�R��e� }#�i�3���~>h�aO���k��A�&[*�F=�������J��6B��7��r��bf��ʠ���й��o�B	x+�P��DX��d�pdGο[��L0��x��id�d��O'�I�a��5��j"s;DzE�)Qw��V�M9�kc�����XH�Ɓ=��1*���)-0��`�������-��挧e���y��+�ܺ�#�-���B��F�?OB+���Q��L0����sF���X$����T����$6��0���99� r~������\�+H�>`k6�@YWk���7ׁ�\UϑQ�d��|�4b9l��q���_��zn#P�4��T�}�@��ʜ���J ���B��o��ҀN��������]}~}��<��60��xY@�_�a�� ��i��6���OG?8��v�oN���H����2��Ǡ������xu�����#@��-$��ghuR�k,��$H)��=����Q��B�<篌x�1����yx���S5���ztp���1�AU�t��^�1m���Y��	Q/B��
���:���:	� ��D��5�;�Z�	�8+%��?-��p�n��kxZ���G_co�&>LO�����G��RI,qk��XҜ��x���ad6|7;��Y�3-�zV�O�%#HY)�Y����3>~
ͺ�h�nD�Yn�� st�A�.m�󕠿���ZM�wdzr�������<����G@+����D1]���Pa
fX���,Q�Z�?�7�:��@���`�\���"�+�������l��Nw���N�2�-ڋ�O�R3�[�A$�C��,J�O���m�����9�l�$o�x_nfI�k¾�+[B���u�U����ڎ�z�z�Q�9�~�t�{����]r���<���倵��0�+.)�W��OO�(�}붆�c����%á��d�G c�d���@�Q%;$<�%zhU� �_q�U�#&�7=���B���� :�A�b��;{�p�/! u>p7��|�o�q�����T�&�Ek�=�U��S������0��R_���f���D���,����,dEk	K��cFԫ岤%x.}73��UeE�5�qS���cx�/adoĥD���w�����������݌��u���B�����򰃬�+�ӽ��f��C�E�}���)q��D�V(*��!k��[e]��L�;�!:7���!w��e�>��Ŏ$�V��-lW��"
\�K���Q�5�к�����'N�(�kC)(�=Pr<j������8�W�[4gH��.�l�nk�ۊ:�q1�f;�2f��������d�/uRrL�����]���(�c[�9�f _��c�?
�L����+���G:�y�ު�n �Ây�g8�@3���r��.�N�b��y����<��Ȟ���0��n~MK�T���m�Ӄ��}��:�e��������0e�x���译?�-��WY��꿡�(�1;`��<�1��l6�g4�e�]�j`&|��Gy���X��3���;�BK\ק�HI硽���3p�5��_ñ�\��Υ����mX�Pbk3h`���5)P�g��v�AB}�K�ze�� �8u��.��.��ˁS9h�
Fv�$T������ȝ5(J�G��9��H�j���̀��<��ܫ0��d�̣*O��LI1u����y`ߧJ>e
�{d����!��v��2�ȠZa����$G��W��F�	�g��w*����2�U�m�i�P�fM��HY��
�]!�R��Ƞi
yW,�ե�_ݢ�c���}c@��g	�S�燅uЗ��59[������{jE�l�B� ���/[�k/�z��I��Ki�ߡ�q�/��%�\�vP��e}~6_e�Б?u��}��KfX-�L�z�z0�r�P,��(C�ہ��N��}�Q$6G19o���. �'f���M����?�1�-�m��Jxd{�[��v`��R�0�7ْ�B��o��5z��R��)
����V�_�Lm�f��liE�u� $��x�����o�#^ߚ,ŝ���%P���=��N(���|�����]5���H~~ኙ�-��٧�
]���`�D�h��Y=M�ƔD�6?��A�y��ƄH"뱵��c��iC��*]��DV/���7Q��;6���ζ�nJ��Kt�@�S���]E�9��[�W�_�P+����s�٥[ypXIR�qB�B�.YG��ɼ����,�3���s���1Y���?򅷓e� �gL	�<�$�C EZ�e�˲��U�W,�1�	i�Ѡ8���"h�%����c'���^OQإƛ�n�К��5h~��4���h#������n��w7]"{��u!Z�VZ��|��%VƏX$q��i<v6�c��c�����G(��5��V p-�à��%��&+���j�<����ǟq߈tP�eq;�dx��,��e�����b��e_((�JKȵ��ٷ���D9���+�ٰ}IOg���=�Ë?0���#?�fԢ�w��e:V���ј;f��� �ry,�\�B�=�	�8na�-�����=Tf�Ū��
_�ކ�������JP���j����b7�.m��ko��7�@,/Z�v���q}����)�-둔��Y��ȶںΌ��+�␩Fk�qC�teo���n�˳p�;����Ȍ��]�w!ͪ/�&L	��Cc��2�F�)�~6��=9�c�'$,9&O+ط�S�۔GꑮCd>���T;���8A�]!?	��`+�ȯ�N��"�?/�z�*z"�T��?�u�-�^�F����
CPKZ��p���^'.
g�y�K*��A�A�gu����k�%�s������!?_�-9'NG	|��j�d	sv5�yqe�y�Бʩ��y[K�䴻f��28��cn�|�[�iw��k��?�>_�ʊ�c��/Y�~�������~�("L��}��R��9/����*�^^ߗ��� �zY]�L�ӓ����f�N�9�f��H���#���1��64�;,�.��t�?��)�GU���Y9 l�Z�'��n�U�|^�������aw�ϻ�s|��
��b��>U��Y��n���O$˒	������}���{����l��?�۶�.�{�0��|�Z�2�������;�N�=��U��ϱ3�pftu}��a����lI$Ѿr�,��49�W�	L>�^���B~������O�ےD9	���ǜ5t�N׌n՜¦�SC��=����!ߧ��'��'z�����Պ�%db�~������a�k����J!�I�v
��zs�#d���p_,ו;c/�~�Lj%�ԅ2$���ò?G[�M	'��5�[P���=x��"e�莇C	������>
W�+�S�|)��l��N7� ���PvV�yl���9�����B'��q�4-QL��������~�#���-�C7�#>}�$��&�����	�dT�{����OO����PQ֒BڸQ���X��:�EH�&JS	������@�!��dêp?�`�����ҕ��T�)�V�-���n\���ABf�lƶD��*J���/Xf�E$m:@S�Wl.��R%c\������MJ�L�	�A�Z�r,���̐�ss�\�W����<,��s���ﾂ�B^"�u�4 �bSV[�vdCb��}AM1dEˬ�:�O��i�Xy��T,G�D:K�U���c�ėRƎ7xVw[[���,Tf��膞�-�^a��fǾ r���{['xoZ�D,jICć���7������Z�l�f���o98"��|�u�ܗv&Sc����������PUA�HI
v@CS�ډRP�|V?f��5Ȭ^�h	c�$��h�;�'��t���ɰ���[�+����m��7�)L�e
A�Ȃ�'j�����e�O3�[��p�Q;��H��r�/�
�<"�&��H����7�����|��L4*���9tfeN�a��`ƭ�Uy&�(�%���B�mV���(9��F�}����O�ATT�YO�����Or���+����Y����ӹ�uUZв������?k�7���̤�7#y �k�t�ܱ����z7�R�i)��R��@��Q?h£.]���+�)_����#A[((���!ڟ����00BϚc49S��pKglË�khBR��4�0z7����[�!EF�~?=\��Շ}����JCTD����Z@��&�JN�a}�@l�|J,92�n#VU�W���_;��5�m�	獇Ֆ�.�Pq�d��½ 6��@	��fO��Y�=,_��Wx����F�}m�� 	�X��iZ����񭩡�D$jg779|�:�}l�m����T�I�S�l��s��mʊR� ^{ݕ���I���eTG��)��i�U�m�G���<~���\F�5!l�le�d��H?"��ͥ'�LhC�Eq�Ÿj�CN�.ڪ�
:"�t��=`�pZ�E# ��6H�M�Ų$��=��N���E*1�cf��m�fu��ǅ���Cj��﯌bpSY��v*����э�gg߭i�g�Ġ[��Ԫ����`���.�K�=�cƗt�[��d�9�(��+cX3����~!s��������er��_������_�U�	�#޳	&È𼭎���I�lJ<�5�I�D���i�֬U��[O��J<�[]-�r/~N*�tX���!��؎��[��ǭ-�/���b�7�~;�X!�U���R���XP$��(�O&9�v��A!
�:���>9\��-d�ɔKٸk�Oܩ�+%1*lY��c����tu{Эh7{=m{�3W�S�>B5��R�{KI\�r��|/���{�������5���꟣����݊���-���ta�[P3��g��B�q�>Z
G�R��6��b�L��yz�r⇃V��sg/��H�eR����Vs�vJ�͟)�x��� ��rV2�?+
��@�B���Ej�1/���h�$y�� 9��8C�ᗤ�}����`zEdMHd��T�0��s�2��1�R�
�<��U$^E��f�Z8�&6��˽� �Y$��M\�~���{tp|��|yn1qq�7i��������mm�}��6������I�O��	�%�Һ�Sb{����o�U��C����*l�8�͖[�H @M.���9�@c�Sѐ�~|�,ԧb3IH�n���>m@�תj��}�ؘi��OAҰ��X	�n��8��L�|�1��@)�U�g0L�+P:��Ν����_>ohyD���:���������G93�:�"��qʷ�w�
KdK:����6��$:��� ʣM�|�5к�;�����	��k������]M`쵴J���grm3�3�ש��m���*H�8�}�Ў=�qT5-R�X�`p�vg�������J6ރ�� M@��E�p�Sc1ƈǌG&�<�C��U�T�xd�l�v�n�5۷##w:�Gw[��Z
��F[�=��g�^<�C�f�U"Qa êĦ�o>t�r`���t虻`����_AYCO*HYڹ��Ҟ��f��EUsP�d��D�0� :!ńL��Jބ0A<�RY�B@��W��w+�P6*�X�)����8J�o�%���Fq��z;j�����J��\��#֡��*��h���]��R9��bs��𥇸z��XhQ3���*��ۑ�⛿��_�ߌ���(�+0���M�.Ԥ�:����6����������76���94t��gh
m=chhA��7=)����n�&�O����Q_ߊ������Km{�4�e1�,�M#`H[�8Ww��7��p� ���c��#�e n��Öİ12�02������3,�V���=E�Y`X��ư������~���b9�%�
?��w=�>������-M��C�>.ј��1,��@��mMט�Rڛ���[�_GW��v���ei�M�r��w	���=i��Y�g"D5����z��G,�rk 7�Zs�zj���:��M����4̬H�2�,��S�x�D�Dc81���!�T0ǟ�l1�����DK�@$�â�X4������ݫ�L��t#�Tbx:�S��Qt���v)��`�`��jN	^1J�[�"6�ßCXʯcxh3	���$�#��%i,'A�<~�0e��M����Rb�2j�n�jf�{;��;����k���T#�����Mt�_H���+|`D߶�'�'�m&�L�Brl�L.���[q��1�:r���E��ʙ��r�$.�9�K����	�c8�s'���1�����:r��/�8�x�����'>��q��$(w}�y �����ؾy=v��Bt��Ns��u��vl݄[6��M�a�uX�|	vm߄m�`�w���iعu=6�.���W�+�a��]����ǚ��v�"f1֭^�Mܞb�kV,����X�` �1gffM���s�b�B,[<K��z�Œ��W=��W���Y�pʊ'�����&�^5E�)�����!�����i��;��'�NqBh㉁��.�D���eBg���	���%��50z���+��5��5`�����y1	
��y�Jt���g3g�����D8zA�.>�e�J�A���b�_ưVP�«�Ѷ�cf�(j&q;C��0 zdy�,�!�ݐ*�zİ1,F�R ��FK�$,�yaɒa��m?U-�a�Hh�zVİ{<��߆[7[y�dAz
���������\dd�����K+�����-,m-aF��������)�ӟ����	M}�SS�����ʱx�*D%�@E��ƶвt�
��i-�h�����-
�Q���񀺎1�l�1������sǱ��N�T�"<>��AP�2�Wpf.�1���c�ya6�62w����L���5�g� bB��L�o6wb2�& 9m<S��tp���3�ٍ%����/_��@�җ� (;F�bxH>��ª�S�v��m�RPT���$���Ň-xɲ���X4��Fmc#Z;����D�뷸p�^qP��a�0	�c�#��>A°qh�r��S���\���-x�҄�G����{�j�f�/ǲ�p�ajZ{�:q4	$-'bڗǵ�a��ے��Ζ���{��@yU5����6k>&��@��jTN��I�+y�.��G��{��4*��G
[e�#nr��aoQ;,�0�W*EB�2Ƨ��
1ʻ�0f!#t
4�{NЌ�1�,Tp}�,��(��=�s�����H�U#�B-�����G�i�Z��PwNA��y�X׊>��/�����c��|�c;6�܆u۾�΃����>怔�;�c�ز[�p��:�e�I���م�����S8qᢔ#g��ԥ+8~�"�>�cg/����R�\��C���kh!�~z�:ڻ��]�a�N���#��p<���F�F^y��9N�n���`�ǈ�f؏�#��0�Q��"W�9}�E3	n{��������Lb����6	� �	�:��Ҡ�7m�0|���߆�g�pg</H ��0W�X�������tuԢ��$�_������(�']��c"�y�M�r���h���u����m7��?n����[x�&��m���t5�`8��z�_)�q<?����r�����y�u��_��+ؿ}�M����&Yʌ�$T�35�aQ3���9��l�?i��İ71AgI]嘇����5�IDp!S���ut)!\��D��͚c���w	a��E�M](�4g�:�!x�>�e�&\%���1� &���,!�Z�#�M�CuOY۰R(��-,�g,Cva%/z�r�:�_8��)X�|)��jP�P�Ä�h��h��t�[���~�~!���G>Ǉ���|.گ��O?��;7o�d�	sS�?�y����J,]0K���jp�r�q1��勰z�BbkV�"+�ò�s����,�?{ �|m��������S1w�T,�cN��\��%b���j~�֍k	�m��
�\���\!ո�^��l	6�^�u��aӆՄ�b�^��7�$��rY��b>^C\�Ö���ݺ����۽��.e�۱�'���Џ�Z�}��cA.�����qA.��j��k�ܷS���}?��3�p�{y5�
1��H��E	�"5n'��ރ#�Yx8{gΜŚ5k��Z�+W���e˱t�R,Y��ۈK��S�PQQA�����!!HKMA\\f�y�9��w�n�����X�l%���akd#=+�����)X�b-&o6lXp4�EW��&�5K%FM'����Y|,@�D�$�	�>'��Ģk(��j�JM%�2�^�a���>ð��p��6����� ��i0���.T,á�B����f��6E%��v�Mؽ�f̚���HTϙ���^^;n�t㜭��a+{kX�Y���Q�{X�"1�5f4�����7_a���Taag[��Ƒ�
cs�PT���#��}a��X�1�C�c���}d�PadEuM������涄��T�U�xX88@��s��Gm�sT�Y%'S���g�\"���"\yЄ�'/1c�h�a��2ץMU((+@US.��KM��9!(&'���]N��?+�q��A�&X�a�%M&�+~��t~â��4f���
T��b(O"����e ���{��<C;/����C�ĉ(��D��TL�(�v��+5M�`X�� ��q�Q�q��u��=1�C��N��s"�b����������+�'��3���}�o����w 6^�P6��ɿb��q��%q*0��C{eC�!����y�4�E������;���=}o������-ڸ���9n"4}3��<���S$+K&��,j������*@+��=�F]��7+��,�b@	�r���ޓ0ƛ`��(�+�
D�ʢ� �*�����{'cl �A�|-�W!Լs0�>YU�u�&`���=���y	��o|N �)�P���M��=GÓ>4�����_�g�Q��ͽ����'4t������G�����=�������W����'>ρ6�F^�껞��I?ں��ԅ������\1�=DX���#���A�;dH��g�����&j��dVq�iʠ'چs;����O��Ͱ�g7�����%��c8_°h3,�V�N�8�P	���Uk����3hik�n���@��Ԍ�!����~N����}��.�Ӎ�n�F1���#��=b@��R���\E̓+RM��Z<�yH��y*����'E<~���%��tޖ" ��~���!���vb����������ѭ�����i�#������S�[��#�����%?��?-�+2�TW�cvi�O��f":6Õ��Kr�����t�:����
vaİ(�M�YX6,"�x�ρid.L��`��͢x�/ ��:���;N����=c�� �i�a;~36i�-Q,���)1_c���	����!B�j9�����V13�0.��0B���;�l;��i�1g�244�������Zbx�ǢۼU�Va׮���C\�v���A[kn߸F��@����\����8�,.����X�>q	[yq�2s1�2�=��N���;��o�>;tW/��{����c�T`���=RN?������k�u�2��gN����p��%<��c��u����|�4n^��3\� �{��۸'���_��e�Jӆ�hk�g�Mu�M�C�=�kA����hn���}����`=:�QWs��?Eݣ{|�C��P狛GEZ�ѮW������.��]�K�{��5�77��9"���}<�}���
���Mp[S���;Z�Yj�Ž;7�=.����X���;��1��ᰴ� ���班[����N��)�013���.��Ma`hcsc����ʱ�'��(����.�@v���{�.�M)Aa�$#��^���W�q��YL�+DY�,$$e���:�з�S�ӧ�3a�g�$�+���D;a�H�Q}�^8z��Y1��~�x�1���(j�Ts,[N�,6�����M%�bx�7	�_����p�4^��x1
��_&�S��,0��*����IBtx�ӳ��w2�R*��91<��=\��	���͆��ƎWWg��z���5ԓ0��� 5�PR3Shii@�����o����̜,�ܽ'Ϝ�d�`Q����
=;h�B�1cͼ���cWj���󖬆��,�(^��H��V��,��f�j���	���5v�;�go��˷a��5�M���X�@Q��Uh7`����.�̹�i�V�ݸKV-�����v�Z,���Th�"5�W��F]s��S(�xq��A��O�Ka3U�B��]+t*���cXj�;$���,C��#�����b5�*f��9%,UE�AGp���N�xNL���g����011�n�stu���GJF:N���kw����/��S���m�a0�,b� 0�!�/��f�3�	а����&p��y�Cj�����hm�j*��m�='��w�Tc;���/Q����I`���(2�q�p�V�yЀ��\Sk�4��ūwq��y�?t7o=@�ӷX��$l#���*aXY�Z���M�z������(��b"\Dd���T�g2�����c='a�W!�1�|��wU�-"���b�����|�h[L���#�|s0��("H���`U!*����=�a�9"�b���X�� �G�����qT�<�y;Ob.�cs6���;�����i�7��z%�f,Gɬ�(��Ӗlƴ�[0m�V)�\�h�J�^��YKQ8wJ�GάH*[�Ĳy��At�x���SR�1<7��c85��H�(z�K�$���1� B��&�aF0�#��,,
����G	���!+�,8hp;�|�ϰ1,��q@1�Kg�]
b^9�?�P��^���J��<�f�?Y��+z%`�KGQR��2�8%ðh���Ԃ����MM�n������~b���^��EZ��YX�}�׍�'��]�?swn�����ES����{�`H�sBx ��W�?�����ǃ�;���0y��|�i�}i�'^@r��~��/���؞��pf�gI�.���%�^��g���?��9V�����v��4��#h(��$ �Ai0� v��LBxL���,�pc�Kb�F�W����\���M���$��4�7�p�F���A�AK��.���#A�#�m�a�^��z�lB`>�"*0R�na9��z'
+�y����k��݋5�8z�4v��W5p���غm��[�3g�����ׯP[S��˗#"$Nv���G�o �|���
o�x��d#0..��H�.Ǚ������Dw?���loËg���߼~wn��C�O R_�H�����c�pc`������&,oݸJ_�5��g���hm���Dg-q{��%	��O����>q�������]8�w��&�q���?u
��ƞ����`�w�G��{��س�{:�۶l��˰m��[�֮�֍뱖�6�5����۰���عmv��^��[6���3�b��u��ؿg7׳[���֭Ɗ���`�l�^����¬�Q�����"TϞ�9����̔����?�cƌ���
��-1!+x�X�n<}��>c���pr�@pX"c0���O���������J��SSq��]}=�uh�gLAQU�,[��e�PY�%��a��S(�6Z&�0v���/���6މ�`�9�EWjC0�?�НcbX4�0���̆i�ǘ�V�,nS��aBXW�GVEO�^�lbx�čvö��a5��0�N�$�Ã��=9܌�ɀ[JL�1�-X�*ڼ����mEq�ԋ���+ƩA�P�nN������LL�`dd@��K��,�`je{BX�XWWz�puvD��/��?��o���	��,��K�-��?��'��]�=r
~QIP�vհ��C1�	��lb����X�z�4��CGp��#4�4����m�h}܉CǏ���f��8�Bhs�3,Z�J��n�t����t��Y4-O^�����X�{� �ӄ�V��_�ݚۨmy�+w.c|N�1��)����#�`*�T0�����m�`U!��\-\~�C�+��, 6�ܡ��D� V�����&����Z �4Q�V��8�4��Q0m>j[;��ҊիV"��-==�^����~<hjř��� s��M�"����P3�����s:좧�d ��k��|XxG ,%s��Ǒ�p��Q�Z��g"s|�p��ml?v���J�Z�9P"8��
�&7o�؃
�D��A�%���X�f�:{���=��s���3�} B�b����p��7�y`��LBC4��mW9�e��xhd7�4��+E�"���e��a%bXY��;�;��`T� .G��<Dw�[<E�s�]��"h:��r��#����q0t���{�]�n�4��H�X�d����}����������|X8�a!%�=kX��߲�=��8EB�5��qR�����z?��J����<�x���Ҡ�-�hxg`�m,���·���hb7^�"�U���[�H7�0,��pJ�Z��`N�o̼�5��<�+�A��G�{�ò�"����&�Èa����~�"�j���3�?-��m�q�q�ax�\�7K>~�4�[�񰦎n&�[i�����_�x!a�y�3�ϟ��O,ԃ�"O��K����������w�,�	���z��<"x���#�w������vޓ�C�X�xh��O���s=��~�5Ѯx �6�5������Y���0�2Օ٘S���e0�$+W#&66��?�Z�M[|�a�a�6e����,�:��X���.*V�Doa��<���9?*֑Y,���!���S���R���9bՂP�H�KƊ�N����?B�Ű���,�z�>ySi$:��%y!LX*7	�sH&NY�̉��NLǒU�a���8q�*��ވ�is�z�V|�� ��X��sb�^B�����v�������)t��ae���{G��+n����O��S(�\�yѝ���6c���9{�O��E��j
*�Tbڌi�Y=KJ���[	

'"R��_�E��P�y�8���s�Tc޼9(+����TU����&�'�}99HNL�FY	Ap�?��=���B��ۇ��A�?�~^��'��">:1QHH�A^~6��dLHCjZ"bc"���_oxy��F��4���;"�C	xy�q}>`�}|-}���8~� ��3�.�pur�����aia
{[��Xq[������f�������4�xy�{����_�����?y��6�DLB2�/Y��k6�'0�:�ur���.�̭������t����ز}7Q��c�1FI��۷����h{փ[��^W�×�a���ؼ�_��������дp�8}hZ��1a,�y%�"��t��I�Uâ;�J��"��W�(1(1,�K���"�5Y��e���\f�45�M-8�����D�n�蒭c��qÿR3,0�J{�c��y!�0�:���"l��-^8�a�HF>@�9�\��{OgG��?�fD����4Ȇ��=�!w8{�"��AOGFz06�Ǘ_�	cǍBeU�����e�������װy�^�:x���t>���1��DmGVo�$�3޺c'.^�����ؙӄ�	\�v�9���Vv�8~�2z_�����@]_�.� C+O)�Z��9���-�=�1�I�ɘ�h*g�7Y]��G���e���������ʈO����x���ų���9TM|�eM�d���13�\	��i�f~�2̊|���O^��|�a��O Xa��R��^���P΅��7�crp��m����߾�
(._Ƅ�,X��=�x����4Ô�}e+o����y0�a�1P5��.1l/0R�<hm<�B�'a���h�iū���uݹm7����ҵ���%�_�FdA�Z�<�ۅ�T T�Es��6�υ�c��?��q�A=������D|�`lf���T��p�,m�C����@?�ۗ��s(��� <Ǣ)��A\<�`y~�aU�`1e�a�DE)��'���7�v�\��;�Lȩ�B�=�Ɇ�G6��8��e,Ls��fC�7p]*Ľ�����	�60�˄����"t̂
`��&!��~�u�V7(��ɰJ��9��!��� 1h
ף�IgA��e5�,(yd`�m�o-c	\ƌ�)�e(�17�a̘FHo�k�G����f�s_�#�ωa���@��L��6�İ?1�C{A�:���o�aY�j2��&R��`Ͱ��h&�V�aQ3���nl&����fx�ϟ�6�����/0�'�?��J���&YZ��^�'Xt�Xs������A����=�xF��Rp��D�@���LO���ǲȗ��Y�`���}�1��2\��p��G��#�'b���U�Egc�و���"@]
�VP4�ŷ�F�e
=+��z��7���p��3O4�a�g"`;��D>O���|���B8%W�1e!:��	�ę0K��?�
f�S`�P5b��Y��,ϯ`X�c~�b�	Ü/B�%΅k�"�{�B�<�A�ḪDRV1\�B��#+WX���y$��������LxD�΅%m5]�H4�CIMj����X����'� �$c��˅W���g��/N�`����M�ED�i�@gw��Y����.���=L�����)�X4FE���`��4��``j*����5�����}CXY[���&�F��İ�����4�� zI9ÇǷ�F@IA�Z�PWՀ*ׯ�8
cGc옑��Ђ��t�-mu�Zp=fP�R���O�5�*PQV�ر���D��!tt�0f�h�5�
㠮��e����GGX[Y��Ó�u l���"^9�[())���6hh��s5���TT����w�ʔ��2���m=}�jhH#�}3b$�	����a|V>V�߂��BrO�֎PTׅ�!��m��	�ذ���s��E9~>�<i�Q������h���X�͟�������G8v�=�ݎ78��y3V@��*�>P�Z�)	���Ãǣi8!,a�(�0\Aˢ\
-��͈X󨩼8M�O\����1^� z�È>�*^�a��>סM��̄��Cp��c��	'�#�aǏk��İ��a�.0�lm�Xh�E@��R5���u,�a�΂�	F6f�
�Ed\L-ͤ�#D[aoB84<~�~������=,����F������pwubp���#!1۶o��c��l�bT�@X^5��E��J��Qn]�p������>�|��mCY��0c�lܾ�Ϟ��7Q�چ��(����O�\�����e�!�:B��ZƎİ4͑�_!a���;$e�������yK�a��8w�.�8�s��`ņU�
@��r�zԌ��]H-�
�P5�a!"
Z�)���"�YP�/ưhs��u�K!�y�iV�D�j�x(�Ec�ԥ�{�M]O��C��Mx��Q�Ԉ���x��\��Ӗ����x'�@�ǉ���e�T;�G;æ���]��WT�J�4���Q�m<}֋��g8y��t������Ö����ʂ]0�$ebG���>Ű�/�����4:vO��������&TM��ЈTM������������_2���*�ݴ!��M�����_Űh*�	����A'P7�a1��$(1���0����-Q4�m��j]X��pZ	m>�
����'b�*q��������J��5Vܬ�s���Z?b2L"�aFԚFJ�����e<�=j^R_��~9,P���s1�3c=2Y0 ��Z�sT��
	ongF�Ǌ�U���X�L��M&b	b�8b��0�[�T|+ ̈�ᑿ��Q��n�a��a�[>ǰ��l?������İlЍ"��X%�]>�����j>�K
�_°�/!XD��x���Qs�����&

����c!�3�`ͦ�X�f퐚�Z"��nA�?�a"X�������~b��i7a܍g�]x�MA�K�b���'-x��Ϻ�_>�CQ���/����C�
��z� t|��ǭ�� ��.2������GR�χ�X�.�������uK�a��IX�x
��.�ʹX0��΄���}�|��W��_�O_��F2���oF��q*�00���#�]`��
+OoXy1�>��񅕟���a��h�%�2"�i�pϜ��p̜��JX�̀M��؈��	Sa�H4�v����VBX�)n��bX�_� �²��DL��9Q3a̓��0h/^a�K�$�c�s7h��ot�wx*b2�	��$�;zCQ��-�����.�1�d{�7(n��p��ApL6��[��B���9z��
����L����;�~�s���_\}�o�s+����>V0�u��nd
+����Qc�kb��8��"u�xb�	���61G��h�Exx4�⒐�����XX�BUU�H1�����줛�&N���Sf`�%HLH����u�7ZC�P���D�䉨�,łs�b�r�����n.��񆇧���c��j���a��(+�@@`�-�`kkk[���crI	�K���֬[�������������Zцw��U��,,[!FY\���p��Ua������8y�*����+���in�T��#��c
sW��X�~;N���k�`��ذi71%��in��ml#�kq�A鹈̫@x�T��Lgf23��-'� &�a%�]������D�f�D����2�b��鰏�>���I�'����&jS,����b"z>y0.�ED��ˤ���£3��ӡ-0��m���7	�0h�A*\��6.�%a�5��ƗI�l��mĀQ�t��=N�>=���b��	�cñz�Z�]4���,�(CWOzz:�o,��Y� e$�fhl k�0����C$�|��	L�^ɂ�!��ӹs�V���S��DQ�t��q ���a�s�D�-������'���	�V��tT͞�B�o��%8t�Z�nES�cL,���L���;Bi���0�t�o�ZR��G7=~���n����4���9Sq��a��z��<�jJ��-N_>��	�\5�mO�]^!�dFk�7EK7:��!�盘Y�'��B��B��S�K0��hp��	4���E�
!p�(q),�ecžh}�W�]�����ճ�������0�����P7w�p+����.l��P�5`�)��5�,��3���`�C��c�ո�т�V���	��g���/����~�g!�x�T8��B����0�:�<V9U�$��&B�{t���}�)���ƃ�&<�m����KW�bǮCRb��[��E��ˆcv��H�4|�F�y�uVJQ��`�Y��2 s_���r���q-�h/�74��$(��c8M(��+��h�����ߩ�C�N�>�]�.�B1�	��8f����p�y��~�1��W	,�Ѫ�/�vN�0�!�N��O֩DU&��7���&�0���@>1�!�XDA���Tr̀��(����B���#
�9)j���x�5æ�0�ɇEh)�R1<B`�T��oM|����6~C0�/���n2��0\D�r���<b��e� �/ ��"Ǭ<C!�{�,_�aE���"�5�Z�aQ3<pݣGu��k@cc�?�a���'x.a��~B�>�n�y��1�u���yݭ��l$�[���nd>b�eO=^�6H8}�~��H���p} -3�59n��&�y��H�!X�X�\6�Y�G���^=���K4�?��7N�ƹ���}w/Fݭ��v� n_8�-�##>�I��NKDfZ2R�����D&�@JNMFVN�t�KRz*�L��dĈ�'#:#EJ�S ��|��$�t��j.�+��*��J`�0ISa��E�4v��a�D>��!!X��D��!X��fDm��R⪥�aE�.AjK���{p�y��9��0s�������="���k�H�8�����~�t'\=C`�
+η��.!m�,��� ��TN,M�/V��p�*�ST>\	b��D8���/2�D�?��ܠo�]+'��ⱑ�;L��n+G�[���:���b|~~8|��ی���P=w>rs���K'hj������K�n������8($:z�0㺔U��G����ذnN=+!V`FK_�`����&/��8|� �'b��E8s�b㠢�Uu�9:@G_��p��	̙���=R�*�`E��ŉ)i�8�s��Ǥ�"�ٰ������:4�oG����"�X��mGy�48t�~K;�i�aبq1V	s.�څVL_�)3���X�a�<���4�E�����Z����+�s�4�]��3�br�\X:����fή��5��y �!��#�'�,���0�0C��d�PX`'jAB���[��83e�K`X�A���8�ƁE��ʁ��x(�$`�Y�c�b� e�xY���x��&f`<	V��K�4:��Ӡ����E�g5�U`V�5>�S�3Y°:Q�[
�ߨ��v��s<l���g�MY���f�z<}Շ���"2��������V�0�����=��03���������q��%,[��H6@zz
�ϯFaaB�>!
&cǡӈ�.g��&^qf�x^�s�"jۻ�`�RdO*���P6�
��X�j��#4�Ŀ��18{����'/\Eg�+l&��-��u�0d����L��
�?���6��'�r�4�_���Û��E��V,����J�p��������{Ǻ.|��}���fɶ���0҈5bf��ɒl�3�'fff&�-3;�����գ�e�Y+��>�M���LOOwOu��)WW=EAU�ʵV$��?��5�v&�m�����!71z0,Z�LY��m#s�l�Y�|�+��$L�>�^�Ć-[x��a���=��N-�khd��9�XFݣ0�!�N��G:����P$o֑<�C���4V�q��YԎh����r2q��Y�e8�u��\[/���-2��J��_>L��CL�j`�ŰUH�ұ����1r�D�5�����x��Wn�/�{��nۋƑ��J*����r0����&Xy�$�;0̈���:n�аjiҍ!�{0��ðh�6�~Z��q.a8�&|�h�PX�؀I�a�H'�<�c�$ي�5Ʌ�.04%áH*�mX
��jxG"��%4N�u�}e1���o5�QB|��D]�c\�0&��V+n�%ˌ���':�F�A>E�㑉���螪���	���0��� �(��1�=T�3,0<�����İ��3��8��؇��=�AN��?�p�n���ԍ��ý������o�x�"�w�n�0��ex��ǰ�_��s�aǞ��)n��|W._C����~]���#H�x�o^<%|�a��S-�_��/���7�;�_=��ǝ�������� R��`U��"�_=��׌7��K�E�|�}]���7�񱈫|M,��r��9�ُ�<�qo�½k��ӳ���]ix� ?=���Gx�y������gp��v\?�]WN��mѺ}/�����s���˸w�����8u�ލ����݇vb�� mg���;�����c���1�}��mfc�4�J	�#�yQֆcB�ӆK])<�����a�ߌ	�!��51����v�b1�qw��E@�T(x�0�� x��N��E�SK�FI�+"	y������ 1lP��3�Y�\Uq���a�T�p���A����OS uZ5��� �dqU�'�C�� ϔ���V�*��U!(6�����'̝�a��ky�<�p �E�n*��@�[���I	ߨd�E9[�0g�:L�������w�o�4�B�$��]<���3������ͼ�ض� ����EKW#>)
� ��Z!T�������a�ոx��u=��u����� <E���~������������!������Yhd$�>>h5Z�j5׹n�&ܾ� W;oa��o�����RKP���@}�pl޹O^����g��_['�Z� %#+�l@M]=��ś����������04�AFn	~غf!��Sf-��·��t��p�qtp��>4�ҍ�ع�6n=�k���µ��m'Y�E�*N��0a�ϴa�άaB��hf��!*}�[����&h̓���>��o��(&�h��H�I�8��L`1���(x^(�P�b:[���2,}3`��JB�3�T�6����  ��IDAT����pOj�=Qm�:���Lh���S�MB�a1.��~)��0�ބ���0P&A��:F��`�[�������� �E�W��eÉ(�k�+��q�F���9nܹ����H����p��IpDGG���
������	���s0~��ݎ;�`��u�0a�X.S���*�:���i���1���F1����z�\�����L&��H�HEYm��Z��=S�3�ڰc��	�X��]��PA��cfvr�ֵ�����z��G����#ܸ/Aa�$'I���29�r	h72�+���ы7p�J2JZ���f.��������9��#`7
����#0,&��fbeN����<8s6�է?a��kP�Ѐ�{v������[����������[K�h��&��Pb�B��"K�C@!��������}T�c�I�|� &͙���$L�>�.�ĺ��wρwH�w`���(1���ҿ�Hc�J-�b��i2[��\U GU�������r��yb��z�
�o�	M|:,m\��
��DX��&��ǡ
�<�1� ��`���a�]��w~?��	"�����b8�ݸ6S7�M��wZ�-�d��o�2@8�Fr��FX�6�*����7�A<��T�k��y+���+�1q�
��G���M3f���.�:t
����P�l&
A�0S�z�D���зC|ˈ�
!��3��p1�rKG?�4p7�%3Y/��|c�w�$>��2�XN Gh1L����̇���ob�)r"��_��A�[���O�C��/<SzF���GA�(�&�gΝ��{�Iq���L�a1��?�a�E♘�VL�+0����o1�����ÛxM�~z����D�B�-�)='��>�����Mƭ����G��ӆxM����e�;^�"^����i_p��]?�ۗ����ß_�]W����|'.�؋�kcݒY8��۱n�������9���6�Il�m��?�s��a��Ϟ>�?|�D�u�P�z�|�\=O����a��5J�ǧ�n�K|$�|S��'}�)�І��}(O �^0�Z �׉�BX�a%_�f������c��|-ur1�+�!,l��<&V��?^1��3`D�F@W��^��U��4ث���	yt\CSx�I��J��EI��y4�Ƴc��f�ed_�D%�fE�
#��1cK�lQH��D�23��iAE�=�H1��������s��s��<���sM 7����wJ��>he>�� �ۺ�,��ȿ����Iwz��˄&�G��R�='��-�BY�ah��_���-if��3��ݤd�ذ� �R���aL�W�t4J�/�V���[
5��x���Cu����v��_)(lڦ����gy�?���UD>G��0�aT�ӧ�Oj*�~)��>��ΟMl稜h���	���黖�t��+�<��i)l�SN�T�d&�K/�9�C�a����Bf�^����=��+Kڈ`��z+Yx���W �ۇ����_ї ��W�xV��Sv�դ�����W��S!���+Y�_4r�S>�p�����TȃC<'�; ���(<�EY"��<HE(X�&�V�{I�EP?�2���)L����F�
YA���gVa��N�͆��V]}H�e��i*�p�3Y����wZz󃫶ζ�8���$�/zd#��RUm��r;%��D��p��&K�\16HV�%��9�xê	3��к�vyZ��Y�w��t��d���_?�i�Z�}W>~A5�p�g;��C����r_�m,���\�'�W���^��[�/����j��<<�������Z@�]m��1DӉf:<<4�|���ElK�������_����B@A?�ؽ��P=�~rJ�οQbz��b�yb�\X���pknל��;W{��G�P��19z�g2@_���E��Ű��.�b�~M|��6l~��և�rd�9�@��LASߋ.J�h�0)��ݩ��?ܩ�|��%M.y�e���)�F��uA_�$����Y�
�V'k���ay�06�|��R�87�����]#�h6�L6X�I�`�m`�)������KDrW�ᝀ�D1��xA��Gb�ql[�c�}��❿cf�����t��V$�!�Cz�M��0|�}�F��$�<!lwK�e�U�\��ϊ�h�~�c�k�'�?����5ן"AD�R�:b��3���n,j�1@�|�ĉ`�KW�����>�qU9R�\�Fپ���E�� ��s��K�5���
ޢ���>���g�'����8r����L?�zg��]o1�蘀W�ePm1ͼ��9>�$��&=
|�����-�B�x�͟��ld�1=SPCx6��۸�O�w��Ś���pߞ��xu���K�'1a�Uׂ������_��/��h#���{�G�fl��,S�����r+�R��:~���W����uő�)�1�@p�,�;�B��(�gi�� Β�)L�rPХ���`^[�T����D�N�8 �[�@7��v��w}����"a���cC ,�1�f 7��s���EQ8^J���P~p���@��
�_1MF����4��I��T0��B� �����[\~H7F0V��>����,�.\g�mkq�1����s�A����w���㌎�0%J{�Tuy���ЗƎ�Ulx���5<Q�g�(B���(������x6Cm�>�	΅��`����R�%DO8�����1N�r^���fg^N?x1PHgl�m~��|��J!��C
4%������IM�����߯i-.��[�q�]#�
ta����F����	ۂ�޸�z�x� ������\�e��_��G��{~[5)	�7ߛ�����'�-���z�vv��0���0o{����>�JR�/9+�9/�}a�֐��G��f����(��7�Π�u�Пr�T�]�g��x
��:���Í:�8�> ^=�>��v	�_��p��']�_*1��x��(���� \0d*����2�A�)o��y3��7%��>�C'�\�p�\����i��
y�i7a�5�J0j�YC��A�Vd�a���D4�3aP����M��M&y���{���t�|�J�
՝\MJ�t{;+Wo�M�5	C%xg2�;�5u��k>͏m�H���KSi�g��@�L��f��h�\�E�b�7���	�֙�E���:q[���_��R�ĳ�pM��4�؇���~�t�
��FR��6	^��['�{��ﯰ��ٵ�fL���.���E�	��aM�o��Sh��#-��Ov�w~J���y��M��[Y��;�0��g#h���E~��zBƙ���p�R�JX�m�Hǐ���L���IW����^AV�`yƙT���'��n�6_���̤��
���u�*�X� ��m�ꕊ�e���'�_��Ԯ4o�	�_;+e��.�� k�r�U�}����:��
�mO�E%22��X�[p�P�=��Z"q?�N�6��F�%� �EMV }�����޿��
�l�db������k|"���^��y�Z��Q�٘��r¥'ʨޤe��\A��*��z[���1I�c���K!	��9���y�2����V�Y��=V�~��=������X�j���|��+����ߔ�%��F�AzQ}M���?���7L�4�W�D��&��wl.��ҙ�ϐ�"��4��*#n� ��+Ӑ�4��)��������1�Y>�i��q}Շ����ɐw�=6��)C�FG�o��&�i�v�G���Sfg��i?@'��G�rC��FSH��>)�^��9_�s��x��a��-R�=)ٶq�Q'at���i��j��Fi����嵎g��ޚ<_�us2�%���ɋ3�Ď���?%([���H~��:���(�w�m���F�e-^�w���/��6Ga��a�� f
^!�ET���+(8|��������U$��sv���(ۗ����*����l�����56�̈́�,���-�KN��=���º�B=n/>����׀`ۼ5^y�������qПv�7A,�B���PIZ��h����%�Ԏ�e9$�
F���$=���v�_;'cB���*qo?�պ�m~�M|�pQZ�\EW�?���"�p�G�Fl�����
��_�ke��4�a����'����c�e;.P�s��Bd��?g�P��<�Y�~PzS;N7#���|�m*�1F��X0c`����6\�c2�6������s���Yr���fO�Uf]��G%��3*!Mz9N?�u��+ү'3m���eXz���
O-Ȥv��(?��m8[y�����J�f��f[���{IAb�H�޶/A���KP�b��ζ��=�8np�0�!��;����m������a�{ �P+��l�����@���6�����>h��2�U�{LY[b���pӼ�V�)�xڋ��_B�f2�^t�&6h�iۤ�O����$��;Ӿ�ˣ�/h�sE5J�MeR�"�8�R�}Z��.!Z0�nZ�����_�&�_�W�(Q9�Y$9���<��$�J�Z	�� h��K�>ĥ���5��DL;�9z�",��f��q�Q`�O�H�6A_��Tga��q���G>8ml�鋟��*��)�Z?��S���ӟ���4�ۀ����D��H�M==gÂ����D���T��e&��g�m��=&P��N�h�@�g}����R�r��5��NԼx ꪀg�7�|�;3�����m�d�ᢍ՝�w���U��x��s���Ӝ�J�E�طXQ(�Y�v�T9y��<�/Y����;^ C9�X=��\X�a�Հ5�,��ͳ����qA-uG���UE6a��J%�5'���>ku�e�j�&
0�"?�%�[�)�10#)%O�[��E�b�w$m��AAI��i���%(Ʌ<��8s1j���l	� 3e���\w��C�UjF����BJpʹO�����+"gTd�����������ԄͿ~h�L����(!7,��>�:�T:-nvRH�t��{�#V;\��O%��g�"��CcU�ܑ�'���ʸ�8���!�e�+n@�h,m���b��R@Y�x"�b*���b,�^��b(H�k6pU�x����'�7�u�DY�Ⱥ�܈{���PB�b��Y�GN+C�o��kn%��`��_9��3���K����l�����:�t�.�Z�z����v��/��r����ob;�N���3�6�7T)yF�پ`.{�|�����J䝺(���A��؉��+�o	��P��S��Å�e��e��=�$𓷧�|e"�Χ��f-��5N�ywdچ��.���,#���2���S�����;�}m�~j*섹S6�����OO�����W�*GMi�K1V��+��?,�H"���Ӓ1pG����f6=i������R��)�ת:#�m�6~�K�,��n3�_��E?Z�2M��q�!ff�F�������L�Tfe2e}>V��U�i׀m��AyS	�pX)��)�j���\C�sB	��#lpS�����_V��:��-�3Scaؚ���Sacj����^U�Z7�%��,�����\�e�/;����֐31�gb~s��{g8u�tC(s��Cv���#��N��WN�ę�E�J��ʮ`��($��Q��i���vI�&�ǧ��E��j���{gA��ء0H��ݬ�y����GV#8�෱f��(���guۄ��i#Z����eBʰ��pmѹ`�+O	���8�A�>E�98٤�qhH����_�ˌg_�e�h��$�r����D� �}"��j�МK��q0����O�fl���'S-ܭ>O�@��;�C>˘J����X�u�Kt�B�5i�3��!g>��O��pW
ଇ��k4���m��]�S䠱� e\X��+p�P�l�%�I���#�V�m� ����ݘQy|��I�zY;�:���7��p�M���!�>��o�����?lz�(=G�}����*?&��W�r���TWU�<f�u|fLf.A�����o.'��5	)�=n�Aa~H�&͏�&1�7/���t�[��S��P�ҭm�V�؃���V�Ū����<�u�KM�\��DS�@�.C������>��{
��c�1���*��΅)%]g�oe�k��(K��ͮ��[���Y�ro�r�`}˂�V~�ej(|�T�f�J��t�jwWL	ĄCpP>+	�_��B�/a�!�%jC7���{;���S��Ro��saS�����A�Pl�zyBF��)YĹJ��.�Sr�Ɲ�,K�D>")�y��mI"�5�֩�v.�ϋ��IIUg�9�wY.���y�qE�[�-� \�h�0?j��:I��Xd������K��u>��N��B��YF^����FZ��bm����M�H�]��~aias��6Շ���2zg��(�'G��Z��R�k,�Ւ͸؞���icA�w;=Aw�Q��	k"*{�}�6���06����CЛ����(4?��� ��Tn�'�4�	W��!j�z�&a��`龧�YD�RV=���He��hg�^l��&�d_��T���A�[��N|��I�hH��N��O6�w��J>������Sg;Ia��*WS�G�u���+e7NrKEj��堨��Uŕ"R���d��Ɇ���5*��D���F�x �{�p����!6v�����,��a���������ö�C�-8&-�����%��Ʀ�Qs9�v�Z����Ñ^�U_L�� �G�4�X�+`�`�,X2��x�����>F�<c>:�~��H���.�Z�p���ݖ���(�ެ\���}Q�?�g�\l�ˏ3�;{
���,�<
��[,״�㍢�;��`���&<����w���ֽJ���j�-�V5%M������:���'y$���^,�d��Bc��Y�c���ǾqQ�%s��.�=A�~���������}zIk�!���l&o)T�ט;>����m_6��5�;O4ä�0{����٧������;eֆ�-]Mɏ��E���w ��$��菶яl�Q�:�V��ǿ���:��Ɠ�๦q�(f�,p��-Yı�Ӯ#���Ot�K��\ߗ�I��71��$ߋ$�
��O���h�w��r+��Jae�g�g��R�]և��`�"Gh�A��s��EHv���(�����]��˛:�?��̊�H |ߟ?lb���"��ْ�A!Ⱥ�����'kw���R��v (X�zt6��	\�%�<9�1Y�$��v
��ߴr� g���4z����G79�ף�/��W��Ĵ��:X���F��`���f�j8G��Z�@>9\* p׸zB"6��E�B7��$M�%N=��ƾ?�FM{��wqx���u:CT��(�g<�d��e"IӶ��;��|
ê �mr���N�`�ߊ:�.2��}sܥ�dxh�qa�G�#����J���EAB��L���4Y��wё۳���^qB�Y#o׻�����w�9��c�?	?��;���l3bqoj����Qʐ�����n8�`4����2&иS���"�hH{�b��i)�0��w�e�.��l����*�os�x^�,v,���"7!�P�z��.���5�?b!����K"}�r;����<+�%��M|oB?�V��=���Ւ�Z\��M�՟-H����<9�BDA"�V?	Q�25�L���d���$(���3�iذWBC�mT/��Y��c�08x�#��}�>�E���m��&'�%���<Hȯ����o��r[����B������Ux��(��N�!��$�"��H�&��j>]�$.�Yۉ�SIM�&�����`�M���& �jf#�2�fN��Ѭ!��4����]k���Rnq7�kzY�+����&��A���_ѓ����V���}��g3��.�G^��14�c=x��R�%7gj}�0M�{�(n6z��it�j����bn	wE�)�6�b&D�Pg�r���]�)jJz���_w�5Rus���Ɩ�����)�yϗ+]8�+�ڲY�ŊH�sO���K�L�;3�W��n�G��2��g�y4{^�c�{M�7�r>1�����[���A9�(řE��r�Ц�V�'H��yu�H^���|��W���E�/%h|�#��`���=�r���<j�U��Q��S�ƻ8�e�/����9\A:>��r�����4�H��cCh�Bs���Y٬���N�Ib��C��K����hU��y�_,E�|�����F
����跽�`�¾'ّd2Ј��Pry� �\>̂O^<C<�u�=�.w��p�<����{���(�Ɇ�z��q���*�6	��4=�8�d���t��-p�z�C���E�C�Ls�(���\�9�!�XW���"5y��G~o���ԩ����2�Ue~Rlvk^B2y{O1`�	���J�P?ӛ����[��Ƃ���>��gBgs��R��L^�����'W�z���h������T&r���	��~�i%��$�wM�=fC]5T0j)�D����S���D�����$UJ��˙R�c���?��`�uJ�`��	�G)�_'��z�	�q�ݬ*�Q~�BR���K�x��l˃
{5=R���d����N��M�;_����Ev^iEF:u��r֤��*���^||y:�Z[�V
��kd�[D�ur���L����k�d_G@x2En�Y��6�I"�&�R��)n���w��|*����N��i�d�2���~�j
oL�x�C��7�2�bo'�5���g�>x�=f�ke.�����Ĥ- P8�+�$��1���H��I.]���Y��0�++�sT�oX��O�����
���f�a�`��h��;i�k�y�˄���@��|A��U��������C$ ��־�d�8�r �]*2@���f���U�p���f_�S���ն�;b�s�`�؍�mv��d�@��h���L��l��߼֕j�=�s܉�^�����S��Y�~.(�n��zm4�P��?�'= *i}��2;$�:9����;���oYL}a���^�Cl���D�]U+�3&��5&�,2�x�
~�:e7��˒aP�ůw��2�;�Sg�G9�*v}l�1�v.�l"��7C�N��#d'w�S�\��Z�A�QG_"Մ�b���?�TT��P�O66��lg��
D�y�rz'��Lh!n'A��1��4�v{L ^���kaR���
�m��X��^��n��pi��YJ:v�ި�)��"����S��
�dv��e ��5?���cg�{�:R�h-c�|�7F��۪N��K�ޝB��7	�"Έ�A`7���4w4�=�������`K۵�C�*�e����{�U�,��F]5��g.�
:-q�g��ʅ[�����Γ��.����U�՘u�kH��sGa��ƞg�{1�ᶫ՝�O�!�q��-|�>疘ܡ�yq�������6v�J���gmw�v�ܤ�-�W�s_�
ݹÒN����)�
��\�l$���3 ���Q��|�/�Emɓ���U�+@�z�S�}[Rr�U���x��oC-On/�ई�)׀����[m<��]�(!(�l�kՐ$|�����%�́D�]c�|��"����G�`=DA��Q�ĸ��q\W1x�s?�v��*�G;o��.����d�p�%얞���y�Ր�>���߱H����_�)��T[�ƕ���T�g�_-�g�(���[w�Rw��rL'�����&B/_��!7� |���2� �_��uH��~`�7�g�)F�&�F�j����@� '`߾U �[�$L>��pTr!�)�����A�{�rS�QQt��� R�b �����p!��O��oc�����e�1p�:��(�JV���0�q��A�T�~�0R5ڍW��U?˪h&��)Z.c���(V�wy��n�3��[9#u�&��.v$)���'p!E׿�u�3Fay:0�'jy"^�h�~��G���T�2
�]"����̉$��s��x5�Y�;�F��Я���V���ByH�-���,�/�H~A�=��T���G�9�[�Kp
*�%[ZC�������&<�Գ� G� �ZJ#>��m^Z�9�,�b������_�r�%s� ���֟���q^��/J$����{���Iþ�+�Uѝ�l�++��9�MOQ@�͓��w�>��ܙY�z)BRw#�Ez1�w��r�:}<W"]��՟��L
�2�Z�*�d����g:���tQ���x̲?hU]n���j>O��^/�=l�����Q�A"r��(h8L��)�2ʚz�Bu�ƿ��������RQ�[S'�kQ�(g��x0e���tf�[�#�]$���R����֚30>�����v�H$R9�P ���f?e"'tb�`i�TҚ�/���	/%�Ӟ	E�ޒ�^�&���S��@*xK5k�����s`����5��*n��o�Ǫ�2�g��"�t�Oot>��F�������.�;��Қ�����-��n�։��6�F�/mD��K�Ӌ�����k�qg������i��@���W��
ƍ�,@��r�Y'k{r"�M^��yXG��-P2$�	��
$ۇ�,1��>3kJb`d(O�j�~C&�g��bfk-IZ�z��0�[bq�U-����*	�;�ߕm��n�8��{n��g6��N�Rt�p��W��7�Z�`��Q4`��&�'xa��H{2f#�!9��@/ �U1��X|�%���!?�sD���
a�HG��e��e���z��@k|�\&��!"�������a����7�a�6�Uxc	��$���XB���+6;=0�i��{n.�4�`�t$�8u;W��C#�}����aZ\1 ��c	[�����y���������9ŸW�/�:?ö�H@�șL������o� �����]Z�c�:� ���QA����/��-����b�*��ԁ����Yr������I���O�~��
��鶺�����w�B~Rvƭ \K�O�L������K�`	�x�}�!?	����V���Bn�\��xb���l����eɅ!9�`_�+�]Tk���c�'_�����>���qVE��{�|;0R>��,� ~O���AO7��v~_�I�Cbv����p�xZ�7�������C�}�%f',@�����D�M?��v����s����b>Lݟ�Ɂ`O�W���G�����~�{��t���#�.���	L��F�?��}�������:�7>ҨK�)�K�4�`3�uap��	�(x�9�δ��M�bT�&�+���5�=��gU�yT�O���مs	��|��T��
��l��������/���Βn|\c��c���s�nb�y�W~1��1oލ��w#��7�섘�A9}K������9 �x�R��m=I�ۤ��5�YƔ"vϫ跾n�5�mh=[�R�����=/� �d�'�	��K���en[^�F�sz�X2��ڞ�;��"گ=�Q�$�V���l���=V��;��ӼyT���(��\ߟ�\.<s�å��� ƛ���	���MH�?��W�� ���0S�J��ۚ O/�#{upk���u���r���X�M�:h��U�'��q��"`�I��+0:���&.�T�	���{i�(���];���lXL�T��b|��@D�x�np?�4���#�z2�qD5�Z{/���P%�����/��`Wy�Cu�r_I;�PH�b�����e�j�ӗ�>h�n+8+��
D2����� L�4���nWИ.W Q�+O�o�p�q��v�q�̂'��qs��Lھ�4�FtZ<�X�G�pR~z wg���sɴ��H.$t�W/iM9�:|�r��5�)�3��>����/ԜU��/z±�`&2�.�n�˻}䟸��99�����ӗ��v�]ڷ�#}��ح����{�(����$��a��)}g\�tzW�7�z�vA�@Z�,���#�#����Ꝡ�vԧ9��M��?1E�?^1�i�337
������TX ��J��חh��v��tm/��TQw�����tU9�{�g�tU�~u�DU)H颌ܱ��90�_�ki�<���B����0$�l�?���5ۑ�ض�0�噙B�\Phj�lAK���;M*Z��u�j��2Y��E�f�"�:l�)t�D�7�$|�f|!8\y�yB�zIN���1Un�[6P��&���<�z��ՠiյ	��2$�+�1cl�z5UynP��{i� �9�͇\�̗^g�����Ȱ�T��c�&�VNҫ�
l\%R�\P�t�Q#K-1�-|�<=tO�/�f5�c�W,��Yw�D��R�'i�1g�m����rM�#�Ma�6#YU���0Sv�h!ģ��`��]8�G�I���9�4��!�q��.u�)�\�ȃ��!�G��8��U��Nf���C�Mz�HR���(]!���o��q0�t��W�=�#>(�A�Y�Q,lRNh�d�."�$�>��9�2jJh%�k�\>[/�K��m���NgF��(ץ.�
���b4Ұ�27X�cts�V�
F�,�)�񟣐CM�}]�Bar�P�ऺ��V��C������g(�HDO�#P"F��Q[���t��]^�ƕ"�'asd2���D�G�/A�S���eˌ%��F&GȪԸN>����!�RL�T�� �0��?��(KZot����>�Q�Bj{B��'�W�q�ӍD�FVtCycyi{�iҩjd�Q�Ւ���K���a����A�H�_mN3���x�~�Q����*��
jX�⥕FS���]�PM��zw�8⣄������ೡ�s��w"��S��l�uJt�P�ܸ�ݳ����]F�n�����X22\����i�h��QlM�+�,!�޼��!�ū�w����7�����Ձ}Ӎ���u- ;����$�<�qp��2L2ۦ���|��aC� �Q�����Ů�����uZ�S���Х��͟���q�R�'h�@���/��]�R3"� �p/1�7�%�p-*���,��C���U�`��l̊~c��u�@x��1��3|�y���HE&�y�eq��R?�]c^?����6��'o�痷z�������Ψ���+��K�OC�	H������5�ѧc_77��m}Zg{3�,J@��0����oܲ�F�_'f�Y��苈t� X�Ѳs����~�M�$ҫ���Z{�x��
�GtX�s�H?T������f9���~����t����:N-Y��=	R�1��CG�K�ȉ@�oє��lNJ����H|�0�4,��B��sa�cA�@GYș���	���M��.�@�wY�;N�E�5�������?���=���bh�}�Me}
ַHE�b���
��L��.H�G���Ӻ7}\qx�"����#:טе�R�r,UWB�c)!ݟ*����{)�۫�Є�*r]7o\��H�/Bc�9�g����V��S�޺�^�j������xh�^�+�������o(ϋ�C�烬G�>�Ζ�;����[x��Ӭ�����r�j$�j
$�(��	�r[oV�PiM7hP�?�� �w�Tغ��f�z�/;���ڍG��"F+�������-=�!
��%�:�k����w�P�X[�9`+�rF(ߨ*�@ 3���|�Z|N_e^]Cf����\�r�l.�a}:IQ��h!��6Ϣ������W�P�apJ��E���<�ڄI�pGk����Cz���j����%$��D��֛
�ŗ8�I�v���D��/I�u�	�Q�M�  *,�3hI�b^ \��/�/�|����B��{g�l�ͨf��=r��[�[&_��,��|%�W�]�o(f>/㖁V��^gN2]���&'ϗ�7�����qc-ln���sX=qOi�6A%���ێ��qt_�fBe���;�-w �s8�A���}$(�U2WVI2y[�݄�KH��TIJ'6a#��RB��wfZ��x��m�,LJ��ܚ1�j7y�w��fBD��ﬖ�	}yt=GcHA�v�,bZ20�(��|�����Z�G!��L:o�������@ԝ�9}��"���,�RpV��2�)m���U1M6��O%Fch�g�EvbL.K����6�s�ci��#����~"�z823��G|8B�"5���� Gf��G��W3�O����$�����g�;���/�b�ZP���<�BցOn-��F9ڸ��2J��2/_�q.Q�X�bJ�'�����^[M)茑D)"�K�U���h�W1��J�dI�s���G�����.=�n���y��:�������\�>��-�hƌ~F��(�����sx=��s<'�JG�ж�R����)���@�W3omE@��^5��xvgz~:\?��2�Nh��M_�&k��v@x�f�V�j-�(�f[�BY8!L�x��H]z~�Z��ǆHĔ��u`�5�,��a�O�n�4_Y&kL��(�{���-j��+�s�ۈ�ɖP�s������2�US98k�LFt9���i�'7��T2��{�#e�	�U~�=qg�2&��d�Pb�%8����Y'��^�!7�$�E�⣋�B�dk�י�O��������ބ7|���Q��)H�vi�1�wU�O�׳=��N�֘�C%� �<��U�;����!'�?|F��<4��~������ș?��4�M�8���R}���G�l�]�T���ﰸ��W�\K*m���������x�5
�����Z<-�AgƖLb�{n��2���/kb������:��NCA�/`g'��M���Yf1&��ϥ#Q9?�o��$�?��ҠR8��p��&��g�,������5a������Q�Y�ѐ�:<H��Ψ��:��LW�T��$������x~}�t(+k�7�fھ���n��E���ñaOEp������J��?<��d���K�W<���3k6�O{�&�AWkW9a,/��ŉL?�~���!��Qi*�}<FLI������q�j�K4����@A�.z�no��j�N^����r*�6�ݳP섀��|՟��Ϋo�ɴv`��'�?��@`��ⓍE	l�ݤ�<���oj��� �l�h�aB/Δ<E����d�0 ����4��\}f�׏͝y�H}#'�ilH���<�$|N��qc˴t�)��K�Y���0�P������ņ}3j�H}�)=S�����,��������U��aմ��r��	���� ��L!&��j]�lh��%ȿԴ���3���.#�n4W�&����y�\�����><�XϢv��^�1�W�B;ŉ������=%�=_���E>�h�䱂�'��'�j�/�&�?b�FCVr����²��B#�lҠ	����Đ^����1�*���b��:��X��h&V���*�sWR��h�a�?��u>,���h{��2���*�2Ϳ��N׶�}l�c�c�5������]�a���=*��BXy��.�c)�ҵ^�7v��ƿ��	/26DR_����D_���(�������"*�ư�W�b���5.��MĻ���1�w�?����p���7C���*EH��.G�˔q"c*�u�P�H�0j?�7ʬ�d�~����x�^�p3[����Տ�({�& |uh֊oct��^^��^�R�#ݣ���;��ؠ�f�of�P��):
�S�?�'0}�;������N�_��=�a�>���J���"�OH�vA� ��p�8���L\�Z�袔N�{���;�&i���M��@%&R(N3�z���IL�c5�+c𚕬J���q��%��] ��Q�� �LX��o��X�I�3�oZd��O��a
6�Ց)��B��n(�<�	TN�Z��Tk}"�(?�@@3{=ꃽ���?�i�P74�p�r�y�E�H�%E�j�td�ILʿx..��+�A�Fn���gƃ��a�.6��kJ���?�/���������ϋh�/�I�jyS?6��\�4�d�0���|��U�]���0�UbN�)LZ	�[z*jx����T��-�")z��O��[�xu�Q|?�v�F�D&�E: 0�g��P������n� D��{l���?�Mh�Y;'�H�����s���~%�~*��WnF% N��g+$d���X2�8��]���1�`�4^��*P�p����7���#���C_��ժ�)�I\����|\�{�ým��K�
������������oo��8��i�B~�Z>?����Sq�Aـ��{<'@���6ƺ(���^��Pڽ�U�Gο�~pCTk�-��u�'�C�:���o�<"]Ka�Mڲ|�*��X^q�g�aOx��rB%��N,S�߃��>п]=cx2i��s6�Hi��i"�Ȋ2č������g,��qR����Y�D�a\��e_�c����WF+"���\�qtr�W	kR���̂C�!l���۩��zD��Ձg���0���L�G��%�.]����uZ��c!]��h��	��婄����պ�@)��x�N��x���<e�n����i
�:�9`9�6������228�ϭ�_'�a��S��x��[-�t�#��j�6e��l��/8��Lq��X=H�hDY`o(P�y�m�d��;�#���XxS>������(���*B���.�r���9�B�;с��*v����v�?�$f��؉�6G���NӋ^�_q]m�:�T!��;�HϺ�Ʌw$A��'��/Q�n[[�n����j5��� �y}6I5��:�v�|b��r�y|���ja�QJ3AK�o���b�����-���ݷ�[�z��e�C�Mɦy�0��" �r�%2:���q>�R��<[�<��˽3�tE��rs������%�&&��]$dā�v缞Rtߝ-�bR^3(7���c�&�������P겫�@�T:�[ʪdt!��3ϡ�����k	4; :�M�==�*�z.�;�MG֡`�n������?��۲�a6�d���8��9����߼�=�U�1sGE�Ce�<��u.�C*���\a��bFn<MJ�ϥ+�L��_f��J��Ib��D\V"i7��׾ZO�������f�oԶ�8��1?x���a��)/M�5#^��w�����W*�EK&�� �;����"�>�ѝTu��Mϼ���,{ד|�.&��=튅����"� �|�5^��f�jZ��Rf�����z}XLS�W���>�	!��&H�}F-	}V��	W�~�(���9����Cύ]\'Ӛ�j��D��N�=�J-�.��`� J@���Y�Y�9��ŔÐC1^��R��'M�}�3��0��WR=<	cer#�&��&�_V,�s`$O��"v�İ*�Ù\V��K�>1�����J� E,죊�*׸JVR��L��Bry�4A�J��`��G闊s�Ǖϱu�Q�۲�_�̅3�ꋐ5�lڄ�׿�u��S���'��t�������d��)��T����|4H�1�m�"�1��D�Yw��r�8X��J(n��g���	���#�����ę;�q���;w	;O_A��%�[b^��I`�!F�Ȗf�3�}bv>w5��ry��f���N���p��i$g����e�8�>�=��&R��	N�, &�H&#ilh��F&L�p���q��~��n�2A����(nd�#�X���/\b����}�H����;��p"\ޡ|��+����/Db�s�ܓY^�x�n �	��Z�5ؘ6!�M4ܗ�&E�h&H[`��0����o�(@�.>Īqo3�����aXw���	�����?�a�����!&���0���M�u�B̛ďF�@�:Z�>D�Of5�;q�_Ge�\�Lð�ɨm����a�����Y�{���'r��W�S"�(�&z�j�-�0a&0,A�1��eX°�0b8_:
�H���ß9��g���°1L��aQ���"�:{f�6��L�,��c8�76W�a1�G�n�bX�/�E�<[���
�����9�^�P���=�p��=w���wvJ�$��n���	^?(��F@�!�)ܫ�ԵԾ�T)�-�{O�J+B�W�`���c��������������8Çw��F�8�{!<+�n� �ͤJ̝\%axɬ&LQ��U�h,�EsUF7ga��aX8�����9��>��%I��D��C�}��P;����3S;|ni����𹩜���&J���gEd�$�"���a��L�'�9p&��Ë�>��0�D��-�
n�Z�DU�)�.ѵ�4���|��:��\'Foh��{�%4����:8ij�F�z���7S���##�!f�#x�[�3�Ĵ�qN�ȗJ3d|�A �B����R���鐩3�G�� $:��L�@LZ"R2���Od,�Ӳ�^^���xEf�Wt�P�b�] \"�NH�Z��ШD��"�R󐐒���\�d壬�	��H�,�W`,ԙ�y'�Ѱ�Eɖ��V�v��pR����CD�!�|��w� ���&~eJ�ǃ�>����J���"��y<�����5���ME!��]���Rd�ՠ������DM�$i���j�5cX}���U���*�V@���5��#2>�E�~�$f!��y�h=����qR
*�0z�+�P�؆���HȫԢ�6��#�	HV�nj����Ǡ��#&LDǤI5e::&�FM�xV��<f�Mcf���S�6)%�ͬgP�r!~k&\I#�ᱰ%���oVo��+��y�9Μ���+q�d'.����]\�t�t���'�y�%���X��V��WH���$�R�����&�G�vc8�D��Κ��[�0����ר
&�Ր'�A�Xg&���Z,<ӵ-ê�rbXܰg��ȘĨJ�aoVT�8�E�E�p</�İ1˰%1l�E���[g4�#���n��h �1%غ�����̜b��`��oq��)�V��^4����뷘8w	;(1��V�0�$���Hqn��#n�1M|�a, ��_���^�0!d��Fp�bP7a>.<x��w2�󁡽�
�0e�,l>��XQ�=w�����"�	?v�=&��\F���=#p��-b�1�F����w���G���7X�e8�����㗠J*�1;��
؅��/�=#&���͹_��L�F�b�"����� #B�_�w���,0L@Yn�$j+�aq�#����x]4�H�ˈ1��}��0�3�Ha�VD��6�x���0lB�æİ	1l��4�wwcX��b���tX�{1�=��B{l����a�m�~�o���ߨw��z��o���g0<(��M3J�Q8!�B$C��H�� %�v�j#���CB~3�ۃS7��H�+��z��S BW�aq����C�M:����@bX�3��c�v4	��[�?e��9뜾D�@^�����ۍa�dГG�z����1��~��p������n����aq����f���nJ���DX�0�t�1Q�����0��W:�1���@��O���C�~*Z���F����~Y;��4�������P�n��aW��M.#��׻�)��{R�h1��\�r���w����"����t���-��C�W�U�9�ڷ?,������q��Q��Ǘc)!�lvf����t4���I�h����̙R�%��c��*t�g"3%V���/>ş��/�����	��o�/�,�>����+>7t���/�Uг��@� ;qR�L�U�Kb��M��,��O<�<�3l���7V��T���;C�+�!0�����`�FdX��!��$֬�,�E�T*�-�9��`��?+|��fx�7���d#�I����*aY7���;Ę���i����GD�/��o�c�-X�n;V�ހe߮�¥�	�u��k6o��ݻ�v�6�=X�}��L�wDB� ��P�@�նc���ضs/6oچ-��c���ػ� ��;�-[�c���8p�0�?�|}��#X�b;R�j`n;f��xx0�w
�_�Ee5�kiC��1n�w�@ۘQ5a&͜��1���H4����VT��@YS
������# ��ȔaX�� �]���'.���;��yg��ƅ�]8w�>�_���g����r�)�q�]'�b/��u��R&a�;,����]��f�f���8s��\��k�p�B'����g/�­;��Յ�̄�߾�{�ޓa��s�`�����-�(��w��������y�n^���p��Y8~�q��w�B��q��k\��'��g�Yuc�i�����11Rf���\�м<��z�g?��/\��c�q��U��u����p��-ܼ�7�>F'����x����tS�Q�^;�hX�%����oR-\�^�-A��کra��r�A|�I��b���<�͊!��Ia�	d+b�B��w�Ñ�e��&��.�I���	���1��N��2�%.-u��'6M�`+�>��\�ef��/Z�!��۩�T�{����{������"�0'����f�C�Y�����lcW?nO,BR`�C�$�̇�'~���&�S>���;	��L),yNYdKa��[��5�q?�CQ6r\�����aejc3g[x�������,�2��u�Ca'n6��5B ����!l��k���k��S'���39}�voŋ��q��i������y{��c�]���5���$�ew�c �]���6�A�XC����9-��qmZk�U��4�W�������x탐>Ӄ�^ ~�:��%�W�8���B����0����|}��σ6�z%���#�#�ō����{Z�5�pa�(A�D�nq?ōm�G�H��5�Mh[T�{ZkA܃�0�E��Rh1l܃a�<���u��؊�#u�u���K2zc�w��{�����0��m\G'R��;~�Lvs�W1�;���WK�ʒ�J.���?��3�1���*̀!�i��0R󷐆��aXD��kDO�D�@�a�O�a'b�^`8V�3��m���g����塟�0Q�m���	��0�A��sO��2vİ#ˉâ��'���t��h�)	����s"��_v�}$􃴡�"X� ��q��q�E��!��!��~"Z��{}��p0�3ZO"��������3��g�+1�D�~D(>f��GR+��_>�ϯ�7O��O�����kR�y��b��_^qY�����3�Y��o_�I<��h)��@}�Rw-�������T��6�G�Ebc�4޹
/����æ�Ӱj�H�o����LLY�E���6,�Z���Yh*#�+�a�w�b̛R����1�)5�d%�ڢ?���_����=�?_����D���F_C2#�-�a)������}`� +yO�P�.�<�`������^qDn��;V�6�)��N��O2�	\7b�= ��48��u7Ty�1b�Bl8���%�2OFSy$�B���yL!���R���mEH�px��B�R�,�^C�	�rBX�z�d�`�KPb)6￀k���Qt�b'Ο>O�î��q��~\�~�,����W�������۟���������*0v�r��^�x�K�N����8u�.�<�������y�2�?fY}��_��_�\8s�
�`a���]<	w�(.��޽�q��5ܸy�7.�ҕ��u�'ӭk8y�(��8�."�񓇸q�&��D�v�_/]MN9��r�"���m�M�D���p�{8z�<�9����#�����s8r�"N߸�;/^��g���Gt��t�c�!��pW�# *�Vo�+�w��#��{[�����6��7b�����X�u+a|�ؾ���N�g �_��7˿���&,G�D�&���gp�a�۸��Ä�c0~�X��0�'M��鳱|�jlٲǭ{�������0
~�È�j�����yF���H�-ǥ�]���1�G�AzzZ�c���e�V&/۰y�6�ߴs,���n�&���\꼋��Q�q��g$����(Z���=/��U�^�/a�̗���a�h)Ά����ڟX&�-�s�����8��t���A�,�	�����Yv��ac0����E��a9��3֞�0�J�EH�ߍa"Ș���S8"�a�8p��ky<|}����f!��8�鳧1�8��,���q�o�F�G2���~��<gE�����Ra��Ǻ0ek�dVt�2��ݐeYL�R�:��^���7���uO�c�� gO���� KG�U�B� &�A�er-Z��(���&���&�0T�����������%�=��g����Ǹ���t�᳗�^����F
<�a�����h6t絅���M�Z3Y&��c�aF�0!D{�o`Xj��kFQ������%�Z��U�HU���d|Nt�ð�&Q����-%EFİCh1L������B!a8���;����Mq�[����u�8&H��&���8�k��z{ �;��a���r��g���C��k}��Cb-�`{���>���0kbČ!���&�Q�ra�m5	��#��9���}@=̔�0pυkD�
�#�x<R�a�E���8�'z���f�G`�P�7\��uXB0��-� 0,f�sND?{b�)�ש"x�>�����Nb��x�7^�pW���^���LC���Cb�!�
N`��tb�a[&��:���I����\��
���x���߆�gf�?���w����E6>QüN�1lAgH^�	û�>O_� 0��&�O�&0���c�~���~��_<%��|.��?��k���������3	�~�&��o��׷D���ӏ��3�0�]��~޻���mC��?����q��A-�w�Ɠ�'q|�*��l�����d�V$`LC�L�����df3&�壑n,K@GC��)ǂ�͘3�c���X䥅��f �|�'|����3`0>믏?�#����s}�l��F6b� GE �����_V�n��g����a
a+f^#Z}c�D�&Í����K���ɝ��U��x�B� 7V��b<]E8�!+:1���
n�b�	� V�\��/�b��$1�D5<4��k�*��D���y�J"X7�t#]7���������a�{�N���ӿA{K�M���S&a��v�=s����+�x+�~�\�q	߼��;���ȌF8f�s#L��-^���۵�ǽi)�V�ʂ<�o�o�N��c��EX�`vnلg����]Ԕ���L�`x�.�p���c�ܹ}�.����K0c�xn�8̞5	s������`���8�o��&:	��?��ū�#.�~�l���;*5#ƣ��S�{��g͂&9	IYH��AZA.Jj0n�t�_����Hn������Ͽ���g(�I�����UL
^��'O�Ű�$��#*2	�����FǘѨ��BUC5���P\U���N��Oo�v�N�:�`d��G`4앁������$2�Sa�d��%ҳ�1�uuH��DZZ:�b㐘��+W�޳�~�4rۉ�Bx��K]C<Dq:+\�@u4�6�	׺n#37����چCL�޸����F�u�?���q�CQE	a���Cwh1�Ű�:A�����C���,�8Ȕ���7,�ab`�U�<g�0%��|���b���p�3Xv�nC}R{0�*C�Uc��
��b��+��R7	e2�=�G�x�%a��e8s���:/�kBpd2ұ��.��|]��n���i��{����'��as�=� ~����?]�L̻Ò���<õE�V��}����?�*/��X�<U�p�����iť(m���*&�1�PFK�d`����wæİ��Ò�[�֕c��=عo'fΙ����b���8z��^����EDrZ�$���w�5I��l,0��u�K-�â���cցP�?�a�� æ�./ZkC+`D���%�sbX��1,����uO�X؏�r�a2@�j6ë�`�x�F~���^!Z���Q�߀��.���0_�XH�����/1N�@��C�X|�J����0'#F�:�><g�����M��,|咈^)DoLx����%s;����0,o�x��ϝ����-=�>��6zcX_�p1\	�^}�ye�S�n;�a�{4lB�I7����҈��j1������}K���ߋ���b8G�aEb�-#�NKLZ���!�w�
�{A����7Љ>��8���5,@�F�'���������ׅWO��ţ;x��6o��x��߹�������S�Ÿw��n\@�͋�}	O�_ǋǷ�Va�������~)�d���o0���|'�g��?����Σ8�}9�.���P_�ڂ	�3G��%���7#0��Me��)��Ȇl̚P�E�����&b���CaV8�������?����~�ӯ����}������W_��D��7���;|Ua�ILCp���!�Bbf.rJ���_���t���d��g$��*I
YP<<���F'U"侑pt��/בV�ڦ1=�k�3�5m�M�GVQZGOG��Y��F�����
�z����{TL�G��2���C$5�3]�xdwhA��n%�J���o<�2+q��ml�q��I�U*�RS�3�`��ɘ?k2fO�IcZ��	A��Ο���`��]���EXV#l�O]1y�*�`��Qp�4���5j
����!!4�Λ͘���k���#'9����]^?
�V
x�B�ᐻ������q��|�nb����팈0ox+��Cvz,�̟�Y��!6Z���*�9s
�r;~ز�Y��d!4�f�R�>׻����쭐3,9�yL>���Cek-&ϝ������8��yN��e��?�B�pH|�mއ�~��-����$��f��דP����e�X"U����5};^=ƞ��a�"�����1L���j�:t ���Cdl0]̈������e�~�wX��2,Y�y9�����&\�w�O�DN�p����àȨ�,�� ��ypꦏ�㿼ą�����d��	�[���W���x����]L�1v��.��ӷ/q��mT6��"���!��U���p��GWL�a�ΓF'1�M#�	B>��ˑZ�u6�XԶ�0�ǐbg��2��50%��������N_���R	òV��k1l�s�LX��Ne��E�ʓ��kB"2�p���z�>v<���F��`��E�{xv>�E��a���Nȇ���y�Z���m���Q�_B�, ]b�ܟ�ɏ�����0��`��u�����#��<�r&^N<7d��X�q��z���C��4��9! nH4bec��1-�İf=s��\��X�������B�&Սuؾo?�^���q3���K	tHV���ANAR˰�Gd7�k�nV��0g�n��?�a-|?:��8� d�����`�9�$	�Nİo
1̤B���uc�Z��J�� �X-��������>��'�����k�m����b�5��^�� p7�EH�����1��n�wG7���Z�aB۷V!�N���w3�T#a����P�Xpf,O���a�o�����ð�����X"Րצ/XN>w�$�c	�^湡�p!�;��^M�z��gv�R7	1y�o1\���m� ƿ����=Qɿ�!a8�������{0,���ƧJbX��I'0�IBzs���I��];�1|��a1]�oXM����߰U�1^>y�珺�.�|z/Xa?t�ޑB`���[�߻&!�܉�8}t7.�<�Kg�©8���ڑ�[qp�&��+����ӸC0?�g_<�)Ut���b���\���N �g4�n����uq�뻃�c��ؿ�[ܺ�Gw���S�n���-�Bke"��(�ʹ#�r^�Ni�ؖ4��`D}.�N�%ߌ��Q5h,�DIn2S��p7�����������``jK;�*\ᦔA��߀@8������nn�
DlR�S�r��P\Y����ǥ#46��x�8��I&��!ce(FiP���+T�@fO2�P�y�PXք�[����Gop��3�<pc�|#�n^����>Ǣ���	�����'8��gL_����&�ˡ�]#j��H����c�Q+D�_�8�Q-�*�(c��߈#�������
7,%,7�^����b��e8st/�ڈ��xX��qm��u˷�Wl.B��է�wL]���cF���Ƃ�H16�\��@_h��w�8�m#�ϙ� ����طc�{��S`o�/��xEA��c�$�ĉ�q��-�Z�QA��N@UE.b�<���qa�3{��Ύֈ�
���g� (�C�Q������ai�1��?������woFL���#� W_w�U`ĔQH�M���%*��p��m��P2r�ʥ��b�˰~�<#�7oي0u0��bd{3�����,{sg`���e���ҕ����7�s�8̝=�o���08���4����Q�>�)���sGue>���R�)S'`ݺ�ػg7*+*��`��#F����}�,r��,t���(%���I3d���`��4s1�g��G~qB�ULBP���U���x�����������UE��/����(�g%��/����p1W!u�S�3�T��a�΅up�	b{"�:0W��+�3����S"Y�% ���b�!9Lވ�A��l|2�%��g`01�]&�'�Y_� &��%�Ŕ�֡���ư�hM����l&�LN�x�6�:�3W/a���ux'��.��mf/ZȲ1sWoĜ5��8�`���v
�r}ݭ��D�EP&��'�u!��ܟ�1L�	XE����R�3{p�I���q�	��{0j�XL��t>x��o�o��wt.��#a�#Zͳ�}3%��=�h��؉Q*B�I��­���ź��3;y��y�4���Sx�3�j�^�B�y��,h�sX�	)ܵ�V&	��ut-�"�6#�M	a&����#1���ah[N{�Q�ZW��\���aH؎]*�C|7�8F|��
*�>�Q?1��"��#R�x=j�or���G�H��!qp/��4ar$aؕ���F��z8�7r��h-��	]c���'^!�������-lE�2x��.�C��<fbx5mh1+�{�(����CC��n�	��А:&-���&\��n������#!��l��Z�"�&N��a1�� 5�ux,��4�<������|-�	Y�H��t�ZL}��6������r�Ek&,��M������b�mTK��S��g��=A�,&�($�ky]�ėÎİ�C��&&� ��=���O�K&��`@��b��8���9��P�:[��.�f�0,Z�����}��
��R�H�G�����-~��o`��\�[�
�����r�"��c�߈�����g��Z�<�#��Ö�p���⅘B��y�/�eh5ᮮ.)t �AX�<׃ᷯ_���gR��+b�/�O���GD����x���4K����ك�xt�:ܾ�[����{x��۹G�oñ�۱����=�m\����K����f�<���w�. �����C��"^>���gL��R��n�#�{�n�{��3|��il\;�([��W�̑�شz&f��D^��sB�\�	�y��H���k�k����	�h�����rLׄ�-�����c����L�Z���1!��+CcK���a�73�p�̛?ÆAF�����G���L�>c&�Ă%s�x�L�=�V|�o�mG�Yˀ�:Aљ�IEr~	*�ڑSUΊ,ުpDħc隍�~�	�=�-;��0z�L�T��\@?��׿r�[���	3q��+\ �KFN�,:~i5�]!���;�������XX�V�5�	A����=�*a�L@r�p8s�v�ELL�4!X�l��oFZ��IC�ϝ����!6�f���k��]X�u7����i"|2�S�}'axܨ�Y[`LsΘ���`D����lF�T�*/r{k���b��p��C���l|��J�[̼&W��E��S��61�p�<DjB�M�V�99Ig8���(+�C`an���P\－_�8~�i�I*CTV!�l���^�b�]�����	�IH�z#���RB����f���t�BE{��u���K��u�V��X�U��]{� 11�	�(.�FvV2�}��tCFj,�3��j	ss=,Z�5��������FN�p%�m�~��B������QHH��x �_��Ҹ���� ���LCCC�9�>�A^h
ZFB�]��
B��4�wR��"Q=qn�~��7����u55�8j��X�p!��u�ƌn�/����~�-�����y���Z�~���qp�FPv3!UKU�C��V Eb5|3X�r[�P;����6��'k�ՠ�;���G+�,ة��"�j#�YI�����.��D`�����0�g���3$0ڄ��pO%.�S`N$��%�I�PMf/X��7����N�=��O�����y~]š3��p��K�p��_P1z��H&��m-nb�Z}�!Z������a��y`6,	X"Y@��7��	h�4;O]��e+�_Q��k��w�ť��p��M�6�܄�����ķ��S� V���Bܼg����t����6o^���{��۵�Y�\��[W��G�õ;�q���M�֊P8�"����[&���%�·�I�o�M�FS��z�k�K-¦�����V	���a��b�������C���t�Ј1~�/�/����$�'`�,z�1�2�OD��bJx=�K$��D����\xvc�-F�J�;�@7q���h�����w��:ĺ�h!Z��k�%p�`]�-ϢuW�-C����9Dw`]3�WLY�:��E|���naq�t#��%��H��"�����Z��C��s;D��b69��8�8V��,����帝�bF��[9����o�נ7���"1,&��%�� ���N���!a؉�<�5�"��/]�a�i��L�0��E���LK�r�/a8��!��<Yp����bؾ�U�%�c8�� &��1�����>���j�e�w�����B�w#X�o�����J �W�.�<0��� .��U���+O�&���T�,{������4�^���a�Nb��M\"�/_�Bw����'�е
�ư�u���b�B��9^=�g�2�za�޻���.����8ud���ľ$�n]�R�@����-=8>vpN�)�ؽ���Î�k�e.�=�{7.H-����b�A������_~䁸{�ۼG�}���p��F��v�t�bXf�c0�.����Iuذb*v���VLǄ�2䦆"%61(�KB^F,⢃�Q�?�|��A��fl۵�wo"��`��%�z�LL�4EE���'�
7�1�娩+a�����gM��}q�`�{�<Z:f�O����\D��:!�Z���A�Y��)�qҋʱu�q\��˿یѓg���A�	��ANI������X�q_Ӡ���;`ˑ�шQ!��z� �Y��?w�f��Z���mPN�P�U��j�G2�eF�TԎ=':�m�a�� ::E�q�HAt���������ؘ�|�@��f&�^��M^q��I�4+�g�
L]�V�9l���0��u0r����P5<� /G{����|�������saf��@x����jb�ӿ��{�b��HH��:""819�Q!Q������Sb�=xy���k�����7M��T#&g8��6L�����eP��@�	CXB8�2㠎U#>;���p��rk�p��U���UcW�7�����d��������رk7rs�Q��XVV���rTU�"7'Ņ�HN���Q�	�����%Av62O8��50N~!�
��Q^4�gc�u`TG0!YƄk��EX�|V�^���amc����:���ܝ����v���;���#��d05p��G٘����훘���ؿ{7�\�����[�N�'&�[X�x&�����!#;7x��v�>��;`� G�8�����d�^)5R�Y1̘��TJ��[�.�@��u��Nc��j�ÖİmP�;���Á��R����8G�"0�M~M�%l�H�0l%�@����zi� 3&|b�l{�p�������3��1y<��5���i�p��mt�|��]O��'�X���@�@��K�ʂ�*[
+>��%�C[HAeJp��2Q_���eM���5�7�>��'Ϟ��Ys��Sy�F�{��\�s!�
��'����<�b����a,?�Xn?ENA�>�X�l	^��$��,X���I���/���Gd#4K�<��!�eX�-.�$ؓ���|r:`� ����R�ƿ�R+�{!Z���^!����F_�"|�}��J���R�=�LL�b*��
��$�s� ���Ű��D̨i♈���{F��;�b	bXty}�ߵ����0R+�f)�����R�V���0, l���J������Ǡ�GB�2, ��"��n�I(��04	���0K-�"����}D����,3������/��$zcXܗ�K>s��6�b�(&d�E���=v�a����EX5�[��>İ��p�q}�V�؆��@�@�DE�	��â/��B� B���v��.'������_��AZ+�ax�h�IFJc���i�c������w�҉��b�&��b�1�
?��ƛW/����x����1|�>�(�;��v���3��2n_?���'�y�$�ݼ ��y��O���;x�����ߗ� �b��w���N�}���kG��N��1����[���]��<��k�`�Ε�yi�^�Mkfb����;+�c�7�X8�	��Uc��fLS�����K��s�:�j�R��ˉ貇���*%�Wa=�a�w���k,"@fΜ��gc按XʿgϚ���cA3��u�HJ� 7?��N���sQZي(B��3
>�D&!$>��#p���پ���
GrA	~�}����g�b������[Զ�C\FbRs1n�<�}�#�u�g%����3����^���Q������U����]°m��۵)-K\4C=sX���\��Z���l?zv�CeM9JJ3QV��Ң84Te`x]��#�'w���,��bʄ�u��n�/a80�Q���Sbxʒ5���?w�}|1��M�U�;ufO��Ʋ2�mnFRXL���-֭ـ+��:f6��|a/�g`��M���'͘�N�$k7|��Ga��:{f~3s|����+���6�6pv��Б�Oq���d6@͊>&w<�
Q��n=��o<FCk:�?S���	�'���`�:o:�G6�+����饹8�uMj�o��V°Wt��J�a�?��;v���K���X����L؃�bك�1���ho����¬ٓ���#�:|Vn
�u��(�}���ơ�q���f�k�f<�'�t?����xqx���b鲕�O$�,m��6��<��S��|X޼Ӫ�H��2�	QB-���	�p��[��z[�l�ݛ7��Q.�8���^>Ĳ9��������
y��u���{hh� ;�JM�I�����+Y�S�T(�*V���j���#�Bj%u T����������9m0�b����51l@�~�6^�V�s����@� C��u	�h��	��xe�D���a�� T���{���\���g8׉���p	N����rZ̦�[�מ�}�E7K�EB
���e�e�S0��;�����p��uT�����m��q��U|3w.��C``���|Ԏcy���O:l�ra�_H�~�9��z0Awӷ����M�=7��Ōof����P3�(��d��L`�"(�.a�҄Fİ�,�N&��L玂cBs7��a* �oİ�;��s��3�r9]4	!j|��S�L���JC`bb%ʄ���f(��	�8�D�+� ����2Q°[D1������v�c�����ږam�wP}���S'�m����a�a��p���uYh�$����i���=�n6!*Es�1�φ��0�.z@��M���-�ZW0�TwC��1L@�����ϯ��q�k�>��d�I���s!Ck!,�	k1, �>�yͱ	/�]T��*��͓0���;��a��-õR˰n������>��E슖_&A�"DB�D��!������ ��_��J��_x��?�DqJ��bR��Ќ����E�a�2|�/�����׵S2�S~���G��ϟ���x�|Ϳ�=���:{�Ο:�
�2Q�PbM��g|��]��iW�4��O�jB�ѽk��y� ���oJ7҉e�Mubt	�����,u���c�J�����=~��`�My����y~�����׎c�wsq��t�:�K��a˺��`FV/�uK�IS2/�ֈi��0�m�su%ɨ(H@f�1��VB�D��Arxy��]f��+�^���Mô���p�|,Y���,ǚ�˰e�:l��=���*Ŗ�k�o�V���-fΚ@D�yx�F�ArzTaI�O-����� '��cf-]��ׯc��h=5#:0�ش��?��k7aβuX��N:}�,�)y�+k����~�:�p�&t>|��rVn����GhnT�2�(Nm�O�((�"��U��Î�b]���.DR�l>x��Ŵi���w��o�
�޺v,�������8�Ɉac����q�f�n=��B�	�����S���_����)Ә���m;p���Ù���o�ft���j�P�1��o���[O�4b�l|ଌ�WP
\�apt���ɳp��&6�؊���l߻�O��c�q��	�8}���ׄ������{�	<}8y��"֢	*��B�w�Cg�/�~�&Ϝ����ș�ض�ej�f�۶��-gB2�,_����ﺁ�<��VJSP+óAt�ݸ�_��Z���l݀s�O���s8��r�.\8�o�/@���C�c��1x��	1s�J?��^�����W-��>q;x�Jʆ�ux�ey�1u"�O����g�����������܋�n4n?z��L�����qy�&z���D-��Jfe��Q�,�m&U'�]��-[��3!�q����[�q��A̛ց��h�"`ll�d&_����+��4r\��a�w��5<~�up�&oe���<(�9y��Q��$V���-��e�]�$*E$A���{����l�Z�E+���>��)��
P�#�kix�X��A�� �g8���m	AĊ���G�M�M�-Z#j�&bS�F��֪j5�RmmEP��(1���?��ys^�������9�u���ټ  K�GU<U��c+wGL��_��ӧ��,�*���r�:�!Y�:��E�p#�?���b�� Y@�YI�V�fPu���F}#�@�o���Տɤ����,��֯_����A��7�ݥ�Nt�V�N��R�A5����'b+���nm2iI_� ����G'���\OT�0�!!&�=�/�j>+K�¥��we�q�X|77_�	3���)b:�������ͨ�jM�rtqߌ��r)[��M��X�W���ГO��hF���b�K��#�[�PW�l^��ϓ���r����R�ޞ�"~e%J��[zP۽V�d�����!
C�S*�sƖ��D�q�c�<�{�뜧�� ����&Ҁ~cD������q��I_:wQ��h7�^��WL����(�w���w!��!�� �Fc6xI%T�C�K�u�	Y��j��$��m_&���O: ����p�.-����$�5��<j��4�=Ӵ�"�q-��������Hߏ��L8!ն��L.ʵ����V����/��(*��U�}�@#�V,��}/���!�O��r�,�t�_z��N���]$}L���*�$���4_-�4��|��"�Hv8$A��e���#�팒ǪC98,cI07L�a0t�~�r��;���R�2��g�n���7QS�������
SY\q��F���4�I���zC	��lrt���E���(�p��#�'�Q�����i%�ݛ'����fp/K%T�3N�.!b?�^$�e���t��� �$��1�Ƈ�W�=�F�;��:�귗Y����$��B�_ym�f9˦�C�6����$��Jh��z����T��'�	��ǔmYÊ��[Apw7�A�-��*V�K�f��w-F&�Y)����L��XG_u(xT���6ءE�O��Eu��b�oG)�^XM� �@��	�Z�O�O���b̈��OsF`n�.��`?l�%%&`�ys�,��
+�P�P�EjVv� 2AZ�&����3Q
�]���H�����5���)�<&�K��~|����!��� �>����l?OV桧�|V0�,��uW%݇r�?#�C�d����-i˼��A.��5�t�h�+<Z�#U��A*q"qLZw�ݞ��@���8JI�l�:��I�jk������nJ:���Ә��+t�0��|xj+���k�����/̮v�D��B�zLkb~&��R�$�'	l�.t"�g$�c�NXφ��/�L^�m6ݽ����N)O�ث��?�~-?�'6���G�#F�#��g�z�Ըo$���e�>[�e2Q��GNJ�����D�,E�j�����������Z ��e��|ծ�X��i�������O�;��1�m6�夘�~�'���>O�b�a����9Ț��T�zUu��w�HNW�Y����W��/'9�RU՝��:�\��ܣ�/��:�D�������Ь"�R�����8�
���o�a3�U6�|��b��5\�G`̡ߥ�ޅrh��ѳr&6Q��q�q��;������,���ˮ�?�����/W2]Y����kj_�P��fD�������\�#zZEOd��mc�8�ަ����}p��|8d���k6�| Q����g<2��>�)�����s�VRM���-ӵ[�F�H���Nه������<���UK5��Ј��Y�� 1��Wo���b_�"I��*�0i�OI��j#0ޯ����E)�O��7ZT���dV��ϙ�F�[��|�~~)�zK/��^U�aN�d��\cS3>d��W/z�����$��I`�A�Z��7��i/�q��z�'Ős��9���0��>��c��nJJڢީۣC9$a͍Lx�c���.`��(��J����$<��~_M[�'c3(����w���7�C�A�w%?��oZ_U�[�
ɥXi��;
aۅRsqK	1���PށRo����(N��b$��|v�ܽ�C�����U 0ȈC�@b�~�?A5$֫h�1�<hL7�M�[��F�t`�A@���}�_�<�Z}���^m{I�&w�bʾ��	����:���q�Z��f�9/68�9�eTe��M�+�tCۯL���5^2f�� H���y(��틏k3e�+�'m����04���}6�ەN};�l�D�7/��Yn8j�đ~��G������ī��RA����Z���L':4pp��$�@��}�2��x��`�6�2�9c�y�o�����^�c��E+z�tg"ۃH2ibR{��HA�YU��	g�6	�q6a!^�\W��T���ͭ��w�f���S�x�~��j�y�6����lJAH��������~��6��Fy4C��<��~��dY9��Ұ����=�����1�#<��l	{��+���ɩ�����-��ow�߄�����w�]�s����e�:8ڸ����� K�p��Yv���,JO˓���npv��"�9��_��ep��ҍ&K��W�^'������q���2���e*��JI�0�C�[ߥ��د�a�=���	G�Y4�{���[�f�-�´-*4�����%Q�rK������������O�#��8s��J4��I�C,~���jaV���9Ɂ�K�UIe�a�@�|�e�*����ac�����{��ܴ��<��W�$`��h�����A WqYX���]k)�e��@y�t�Y vA�֩�1�e\V?;��7��3X����I�ΧG4���b�E�'D4��)�����w�`ׂ����0[�Ҏ�D����h�3��e���48�7a���y����?\�K�w�+=���� Ҿ�w�z�r�������*5fg�mԤ�T��g4K9;�>��,yF_m�����̍m<��[�������ҷ^$g�=�IZN^��~2d�Z�����H���a�D���nY|�*~����{�,����(��B]2�$�����_��>H�J�W@��V�QQ��'GtZ���T\�=����4H�-�_���U�ū��A~��&����2��k���C`^�=�-��~<��-����E��pa����/��=���x���6���#�2����_�I�d"6�q
xl�+��4�Gl=N�jrL+����j46��պ��r�I"(	?�ny�t��Z�p�)�\b�����r'ˍ���)v��� �cm� Δԓ�5oj�ʍ�&�V����/Yա-aS�:� �2r���IJ�X��r30���Ӡ�܊ح��j����9hlS�&�z�b�-	�qT�|Ω�� ��\��S��r���X���m�k��NG?�K�6w&��t�%,�s��ȿ�@�,i�R�����+�8��Ƙ῾�v�h>�Hy``�\�O�ij�E��wh�>�潚O��G��T�6�`Ĺ[f�)�ʛ�Ľ��3�`3�
�q7l�D���SĒlfo{�5�A�iϟ�[`E�гI+g��P�烥�a���^E�"�w�w��r��o������#�(����Վ�����5Xň�p����]���#�`[�&9����}�q���9�� ����V��d6�b�"�Ƌ�He*'�]��0O�$�r����叀�j��hl!���|��}�s�lͪԾ��������s��>��|j�'���7�=
��?��׾㶲̗����3,
�Wj�����A�ȣ;�����~�0m�W���������׽��/�6&�2n�F�Ҁ�>�ȩ���Glz2y�6�����^�T �����c\�+�ɳ����|F�:���"`��]m8�Ӏf�����;��jcq���6�0��N5�i���h����o��>xU��{O�pv���S����h�U�#�
*�\)UTظ���-�7,�,(���&��(a���;?8�$�V>y^@��~�J��FA�M��V<'�c#����xd��z=z�Y�͸���:S�{#�ز�8DK����_��gT�dhY�k�����'֤"�^�����v���Wd6qc�vR���)fC�a�o����h�W�NlP�h��Ig�A��g	5�Fo$?�S�{?`����'U!��p�ؖ���{�J��bE��&��Qʵ"3�7ic=���D��^Gŀ��d
����!������.xl�˳���z��@���/�~Y��q�tת����W	�`���T�%�0;�E�ݩ[m.}�4#��픹��uD�����:ϴ�u��}���`\�J�P�����\��a��||XJS�Md`�փ*n^y��t�?�<q���������sM�`�Ťx�3�����t��a_����3~�~��R��}ʞ�tm�i�h�w��Ή�T����f����fw{$��1���$ç�udc��9��B�m�{^ۚe���stJ+0�z���U0Gg �"�䧶 C���ع0�zy6ܢ�h��cl;��A�N���D�H���岼���e����j��z��D9��*ֈ�O���]�Acz�Ox���p��u��A�H?��tt/ɡ��x�U�����?�:/�y�5�>��M^·8H.�K�H�n�|0��=s{����������b��!�I�il�!�K�\l�+�*bP�Qػ~���l�4� 	��^{��J���m}�/��Z��l4f��]�#��C]�C-VD;�����t��/	������o�Fw�uA�"��˩��ҫ-��}_sq�yݥ`g�S�g	�QN0�V�,z���x�sa�Saѿ�"��)i]��?���M�/Psk�*��#d�k�3��g�Yf�Ӥz�R�jfלܨO��,�
q�����b�_��
Ir�i��EplN��~�@��'�o��eS�8�(Ѯ�k�j~�]X��)/�0_֑�m ��b{�Dח�l����W5o��	w�R��[�tE�cׁ��?�q�} 
� ��/�����.�b(�@�ōw�d�2CDO#�:�Vt%S<��1��w�nЕ;���R�nE��c�G��eh@kL oGJ<V,|���A�荠y0 �_��%}��!9{�_�W�a�sB0���,Y�{{�\Щb��>_�Sg���s������/S�0~�eǡo8��D�݆ٗ��_�b�E�������G?ǨC�>uQz]s����3~��_QȨP�))b'&��·�T	�`Mc���΄H��_~�~yP��d���$SF~�ő���K����������3�f�E��*��:9��|��{x���<!���������v��r�Ri�8����U5"e�W��^���y�5�=}B�֏g���2�13�i�w�ZD�a�珴d�Ӱl�;.Q�����*��j�(9tâ78�Ԍ�$Vi�(�P�DB7�+^� �~o�y\�Y��>0�_�;�|*���*E^$����g�p�$ױA3v�AbD��ݴ�x�j�w�N��3�l����.�F�1ۆ�~��q"��#ޯ°��|!�2J��I���6�X�̮��4�	���?4u�b��e?c;;�R�b��#BH����loH�Փ��JYQh�J!�D�(��4!��2�'��ٿ�O��"ڻY@8�d[c��%Ӷ�k�)�EȽtL�Z�^)L��r����xN���[?#��"�����5�(�z�\�>��c��v���9�>��׬M���Ÿ�(���&����h!�5�|�Tw���	K�5A������Ķ| ��膧�[�����;lt�c��o��F����+�����G@�3����8���J�F�s=o�@M�,ۓ�?as�'�3u�Ac[��F��hĶ{��D�gű3AƇ4�1�!�6k���W��
�c+��fq ��<����� M�Z�h�o�pkt5f6���:�"�$��X�Gi�3���4:�F�ZU��u?c���@P�����)���zc�� j�qa4�J�!�y�4@�����J3����o=Hc���wK|W�����ܮ#����kݟK5L@��ܡ�7;L6���fWS���	�״zN�'Hf�I�>���.�|ʊ��0�ע��/�ފ�CY��H����>9��#�����թÃ�6���$Q�Ŝ��;P���<<��d�4�`�:��/������m��B�7W%�ʷU��{�z��0��v��y�*�Zj4)�d��0�~h5�ܲྶ�۪n��d��%^�q�@�c��]f�����f6�K�ND ɇ��&ۻ��X�\��wa��PY8x-��Yy���t3UUl lj���u��:�����
��åȩH�^X�7/�~xq����f��=��!64�����Yϙ�������S����z����:���O��/A�<�*���Fi����}��q,5���,H���c�3��\~����j�Fܧp���w�%���Q6�����z.�;"b�OIѭrnv�b]�ZM�K���ܨ��g�x�H��%�a'�S�o���%���b��� *Z]/`�dQ&���U5�}قc_�#d��ܲ�HH^�R&�I�r��cN�G��-��ag��ԥS�<O8��Y��8�����3�f�&�3k��2�_iG�Њ�!�����GS�8�@U�����N��\������2"��8�-��9��Ӯ�����T]bS>|�=-�\����w8�z�Ӆ|��5M���]�E1��A)�0Mↆ8��mEa/�\�X˫~C�o�pp�@�QBR~����S��*bc�cM�`M�<�5+�O{�84����{껍)��8jh䟈�X��<�[&�|�/�L	/�^��Q!Xx̿�v��Q}X~�M�g������A(�S��N�zhS�����~)��z�����m� 2	ԣF����Xc���u<4/nx���"��E���һU����_��6��4��+�4
��Dͩcg%G`L�)N�^|�,�"�I��D�甓�B;�~�:&�IM�_H��xXN;/,�G�� �!�<�L:&Y�6;Vӻ�������l�2����K�Um�DE��#�b����� _����^6�����P�~��ʰ))��t����$7M��Ͳg}��D�Xb���LP���?��\<�֣�l�&����Y�	T���O�S����tJ{ҡ.g*w]�]V���$���Q��nf��V�}��\�Sr����Ys���N�2CKI�5�A�s~ �O�ނ���h�}EA���`�s"���B����gc�v	�w �l�}3�S4bN���!��*i9:���v���t�p8DXC��&�C�Ӌ��O!��1�A>b��FND�����x^�0&L��=��S:qw���ƴw:O@t�a�h/�ǑZBM��50�/�<�@��G)�n��&�O�p7�WI�=�C��.����t�I�S��w�a1�Q�se���ZP���(+�і��MG�0�P�R��-C��`)�JgK���������Q�� \ �3	�#Ɔ(L�E�u���E\�ݗ�e>y˛B�䞂{�r������h���t��F�1���y���\�v�32����H$34�VT
�	�<l|�)_��q� =X�#��������ҟ��ww�V��������]S �eb��s���)Š?�jK��_�{�I,M�M�����qU� �5ًhœ��(I���=9}Y�į����Mc��}B���^õ��ѽ+OiE���VZprt�S\&����������C,8B�E��8�|���I��r���~,6��o>�sOE����1�cjUL���#�)$�!�8�������i�q��~	�Sx��s
~%	N\��e3uN)D����"MD����]�R�h����U��<��m�Pazɓ�>�F��=-�ozڃ���W��%�w$D��Ť8L���%��98�:1nl�j��"�N�t�rx�/�����%���Q�k�f�>��BJ��л٪㎰T��d������<|��i�P��(�<2=jYdc&
��}`�p.M]����c<��	�4Ì?������������ܥ������eb��騱�&��:Z�9��C	R���[��a���3�����-?�u�A�
���!���^L@� ��X@R����ؖhh��YEp�!�49&�OQ�}ij�)�ܮ�	���T/�
��҅'>UHZ���״�;v	˼�{x��'ipP� �4�}H��܎�2m���6�����Di��<��8V�'ґ:���n��(���%G���JRN1�W��Q��I&�ZHG�.��x��t]�)��݇ {X�x<��o-%/F��\Ѐ	����v�=�@�|��FQ�RB���*L #���%��H3�-m�ͼ��ˢ]�.l	��F�x��y�	h>6�W��Q`�t5f���|��l��X�~�󄣎?Q����k65��^@QS?ʣ�٨z�ua�Η��*�@ὃT����F7Jo3dۻ�v���(�6�����j�L�w���^M�a�����{c)z��&������XM�rbd ��g����x%u�zkb_�O��ڽ� �8�Aj�C�N%�;g��s���&�H_O��U����i�=�Y|b+F���y��/w�~�9���H�=��%6����_!��K�ב��d^�l39��4�j���6�/���{�>y�Mc��z
IT��M6#�q�..#�a꥾���yKf<�0��M�r��g�Gt��?�JP}��s����߳c�^&��^�u��s����76�8��9#qZ���S�D�\�X�}�J��ܰY��Kfo��hyW��}��X�g,�іf�_��EE2�ߗ��4��������)�oS����v]8�n���ot+Z�O�5Yף7������yˑ����'^��f�f���{ ,�9��$Ϊ?��s,	���nb?��K�J05��m:
���`4�(T�C�uｵ�Q����g�_�%�}(����l/j�|�D�k��+�q�)Ɵ{r��	�菌�I�VFnq��p�_��I�2I�A�?A��O�bY���R��	4��F�����j��h���ѩ�_�@��c�"��	j�B�@��v �HF��'���p�暃%Ֆ�U$�h�}�iy;�Z��8�V��LX;��'��ῤ~��yr儇8]V�	�s�a���+o՗hp%��(��<�M��l��ۻ
:tt5�����dR��Ј!�]Vey�o�]S�I7}f4���q����Z1�u}�L��@��q�iؓGr���Sc��|�p5�th:B{q��lRʱ��d�>ex���㍷�� !��(��([T��W�	�N(4���ϵ����h�Ħ8`֠�w�	*Fn�P��N5ǠdY�Aئ�O�P��vA7�n�x�tE�	�Y[�3��0Jah�bT����Ʃ�w�W:<�`#�dg��!
���'8b�����VZ��1>Fa�'8*�P��AB�_����-qVX��O{���n�0�cD���x����Q���ȸ��7������씦5���4�E�l�=?L����I��Ư�.����U}� � �;���O~��P�_��W�+��Z���pĿ��&.'UF�gw�Bc�s����_,[�� �4�jLW0�Y�����}�e��^�����IZ�"I�4��O�gH�L�QV�v����e���W �[��K�>9h�lZI$��VlYvDs��G5�u���O�Ӯ���}�`Tq5q�� �M6�$��;HډѶ-�:xk���OI�5�z:)3CР�����uu�;-���n���*=6)���*|Z`��@;= �jV��x�U����C�?�!PV�TV~1X�4�Xe�S��;�B�m��۾w��Zw#�5�v�������#i@��8XC��|4i_�e,�0��$ 
��	�)�KB�b�P7�ᕩ�n��}h��!�X�$�;���Ck�KӋ}D�O��2�ڜr�!33�r�l��}sj&��Fn�hKv,F.߁>I7[���C��5�XT6��cO_�P�D��lK�Vf�&�/{��6;j\���Z���4b-���bݑ�mRV�?���,�w"X�6���T��h��9`0.�$?�C�3���ݛ�u�А�w�}ማ{%�����!oćl٦ �|O���{�w�'̣`BwmDt ΰ���^��k�x�/?�V� z��߽l2X��Ӏ>�O�\8s���R�^SqdNXT;�A���6d����Tt�&OtO��:h)�'��>w���D�1���I}����ЇQ�R�}O��o�0�5g�W�fB{��a�t��WKO5���`�!&�ie;F롕2jg��W�I�޲8���fG���,�-�uMzw�I���Q��΋��^|�����4>��-Y.���~,O@�-��|.�+��,��$��h�?PB(r�>�4{w�5��ۜ~V0<����w�y���s��"I.���bl���0�>�2�AՌF��=ڇ_νB�݀D'Pe$���1��5�3���W����~��Z2��=��-1�n �͖�O�¶��@��CҹLAw��u֛�.�_0zҩ�֢6y������{�w�aA�����Ti	�E����V�����{���=�2D��B�i~?},Ԁ�;��ݺ,"T!#�¿-�{>�w��L:5&�;���'Hgpm��b�?�(����:1L��D�����<C��hKe9��3��h�Ǆ+~}�5���s�`��;��h��W/�K=�˶��vCo��9��1v3��Hǧ��)�(�Fts�E��$��V�^,OȖ��s̈́VN���2D�4�b{nK��5�ސ������W&��)���]+`�h���,��$:�{���Uw���,�;�ީ����G�#�kJo	�:�ӆ�3��k9[w��D�V�s��}"��y�@T���Y�{AhL��N�>d�Y�HP��6*D�QI4����{��!���#I<e�Bi]2pq�߹�Z�F~(9��Lr6.�d+���ϙ(�`ea�&�}?�!�=�d�4��`�h֎���_ �׎���W���>r��T!�ؤ$~�����r6l��:me�i�O'��H��z���A�_�!�H�=5��bF��������=o�f�{SW �Ʒ)Q�:8�|Ni�G��Mw ������_UX��*ʂ�v&�  �u���d(]�=`����S@j�FP��ڷw��ߕ_u���u�3�N�S��]�^�"�(w�� g{C��#
$���Etqu5���ʈp����9 1��(}T��2ĺ���͛��L",��H2S�ƺy���ք��Q�D����6�3��.�����������_/]7Л�� ��n�{�����34���e@:�P���Cʐ��{�]�����OLɆ��+p0�����'�ʌ�Lb����70
8�˃)��M����:�������=�X���8[��[B�ƂhL4i �'ǭ���>�s�j��Q|5,@��GEQ���Fм��r'
0��X1�#�>��&O��݁-fb��F�c�0���`�d<ѫ/A�Z�4�]O4�~��q��ҋ�<�Zo�b��P�q�%JљB�{^�e��w, ='�����n�df����I��O�|�
�L
�#��Tu)��P�l��&�:%H��P��o���je��g.��ݻ#�'{|�%tt�:������K!�(���Ie�5w�:Q������#.���!tƫ9M͢��7�k�x l�[���_V<s�.Q9Qd�=����X��l�)�?.�+��ݛ˧x*ȉ�=X�o��sF)��"�]QNX�j�Ié�sI�	U���e������ 6�z��16 K����e�����E��x�<OO
�Q�ˍ���{.�۝,M��T�9=�w�eg�qXL͊qS�ZSe���*C�~У��𐻇�w�v�:Cm�Lڭ4�ZLxl_�0C+deE�/D���� �~�UA����_�Y�@���D8����z:�{�1��܀T?[���u���>8��T'�{�)$��$ �-%�C��jh�_@�����@��s���<��5�X��Y/���-z���xj�9��Ha��,
�����wˍ�� ��$� F�tF����Con���k���Rb	�-�wxO��0y�2�h{Yº�BM�p�&��gg0�7�p.V���@��}�@�=�,u�w0�R��7��������H+�s���R��B�s��Mj��<Gm&��c�=>G� �G9~��t�yŴS�	��Ͱ�s�}��/7�����kT?��I�?��`7�7�2T�Kz9�M5�#EO��@��%>�)����?D�U��̛��k�2�:�39;��^�E�D�?��|AO���!���B�����.s�.M���A�s�LW��:m1�!M���4��E��orL�S����������{l1g���~�	�2]|�<��r;�g;��^�.���KW6�wmgG��%��	�m��@_���r���P�z����v4gO�Z;ǻ�ah96�e��f��լ��{�xY -@����g��zy�*"�Vf=B���8�^�I�1��YF�ܶw���$y�*A�j����p*3�rG���Tp�X��7��+wmj�{Fٙcr�+��-�\xB�h�8��>J�/|73�P�J؛��_��i0#k�	?;�O�{N+|�t�bL1�Z��pދ�S
�]� I�{ǫ0fx��Ζ,b9���q�$�:�u݂^�����g�.B��=��S�}Ʉ���nKgs�	I��t�]&c	El���j�u\��,�^k=7U�wI{$�������¥���_�6t��CA�PЧ��#���ܴ����<kl%	*���N�;�x��1��(�Ǌ��� v�Gk���;<a��Y��;w������-������������ô�8�p��m�'ϩ��O��~��������˚�T���U�#�Ow1�z�<�����Dx�@S�7T�qQ��5��j4�4�$���`��� �d�t��������X�XD��g�^���L���ܒ��'��%�̺��B����Bp��;T�@�ǁb�^7�_C.YH�6�t���%_0~�Km���Bt��:�cvӈӘ������}x
/x���u�e�2$�Ɵ�k�S+ˊ�)�11�!���R�H,�8S�]m�fz��ǹ���L@��Ϝ����J�¢�Z1�O���I�}�B�v����Y��SL�Ty_6�Sf����K�w��'e�8�zf=z&F��,������H���,s9��oJ+-)���ǜ�z����ndr�sR��!ќ���HZ��a%D�,��S~�t5o�gN�^<��^��Ջm�?.�����x`��X���E���Zq�KQ1b����l+����J�W@I3-����O6x!��F${>�<O`�]C ����I@ܔ��(����	���j���^�kP�>a�N�������Y��k4C� .&�����h��Q���"�ps�X���Z��\4;H̫IĠ�j"��w������������W|ǽ�D�mK�(�֋��h�N��	t�[3�уŽ
��PE5��?k�_�n�W�*!Ͼb��6�<�bG��篼�}Kю}�y�T�A`L�g)�o�2:�$��>����"{z.��ɉ<M���^8;J$çm�8�D���;�l�	�,�Z1�_',�G��F�gS�Ԋ!��{C��T��^>�
=P���"o�VI��\�VK�)�/�#�Oe�./-���u+5Q��-�d�������XD"Wl"�C>~c��I�q������MALg��Cg�~d��"O��]zb�B�(>ݓ1��f����f�=�K�KQ�̈́�ͺ�����Vm�+֙��-��0������~ �$����/V�*U�W��:��:��~=��$~|'�&Gi9�j*�Q����1�ӊ�49\֠�
��up��U&�s����`�}6"��
���M,|O���Ϙt��%��
�Ǿ�~a2�`P7_hO�٫w�]^��.K;�:Υ����E
AU09� ����AtR�f&r$ٯ�Fs��{Od�.�O_�'�˻/�q��SEi���V>�"��e����"��;+��5|b[���A����fZ����]	�cWtwd �;���B���DUߛ���F���2,�e$�nw��ep3�͟.��D,oC�}嬮h�X
�}TSh�
�`{6�N_���W�=����x�Lm��a�񡃅�����j���E4���̂��?)t�%y�qx� 65��+����8�)� �>�#���[�H�����G�= P@�����2�3��S���%�E���J2�<ȝm~��L�K�>	u�L��`�)]���u���P���&�&�����e�-�r�/s�:쮺gx���K���'y�9#�72�K���r��&'<w;mb�'�/F67m�C�_d��(Z��'�t���Iܣ�Mx4�裠�3�`�=�[j �GC�tJ�XO��s���2Am¥#�H��6��~��xy	(��dp�i*1�#���П?Ӑē6��E��Q�/�nxK�E�8�W�s�����mwVj�@��k�2A3v��9��?�= O���}s��%x����ճ�ϥ-���5V�{�+|�RдU�5qcK���LV��6Ol���q8�oZ���
bg |��:�Z��y␻+����h��E���[�$�e��ɓ�}E(�Q�H&.^��jf���mJt��������t`m��{��B?����B;(=!YppM�f���/Ȣ���W++�PЊ�nP͕��nTs�����(T3q�t�l�h��4dDO�Cf �e�;���_)���[=�+�	����[u��iT$�$ܮ����r�Л�g�aG��4 �U(Xd�� ���T�& ͼcm�J�Ӷj�鲰Z��S{m��EC�J�A�ք����q�]�s��F���1Rl1��;�c�����d�.�V?^���hH=V��z�KxӼ�&(�;ݛ�ցʧTU���7����"EwR�����Jۨ��q��7��az�ђa"7������;�`�2k�r/�P9#�"���v�T�y�U�.�+��>t�|+\����ʯ9-
��pm��bh�[�h`K
e�hmB��}�)5��|D�c�a�
�bH\��ۂ�4�G�X����y�)]��V�/:$��`KCR��s���>V�|��2P{��h�����!Y<4��`a�lᄡ|����K��9جD���2�=���y'�@[�ց��Q�`�*10ū�����ql)�)▪X�=� X$�5f�X1u�ٰ��b�v�������s�~��:��l�P�/�����O(J����Y�r�_��������ۼ���j�&ϟ؊�Ow�	������$G��6m �^p���W�J��v�h)Pn�
C�/˲W����\!=W��ک2�i�"|I�+aԤW��=j��o{� P�	>^�i��,q�^vc�G��3���Yo@��?�<9V��/.�OT���	�"��(��n�m�+֘���%DV	>�vֲc�K�XY�{�^ퟤ-E�h�[�H;��!aI��I��F0������²��)�*�fDM�P��^ܥY��>��[����\�O8�Z/K"&�(�M(��^e�]:u��j�ǯˎ��a�]���^�R|H�����dɽ��7=S
�d2�uC�.}������UÊi\r\=��P�9��7�i�r����Y%/)CX��X�iJ8/�s6���l�d��ߘg�UԢ�Iy��A���+peU������ G��Vb���lm�8�%+7�[���>��g��:&g ����p�~�`1v/��q!V��E꾱U�i"��(��L+V$a
�5,&ҋ��a�4���7�,��N��]�����ؑ��`�8Smݻ$�x4@������ynjF�[掦hM
�Y1`Z[t��$�?!Yk���D����nG�̖1�b��Fԑ�����Y��2���1c��K��绸�����Ϛ[B�����M�2�o�$�A�:I��@�M2.�LY�'�w�?!O��;�IK�R�����<(�&̐W�JK�g7}���,�������I6�<��d��eꯐ��`"!���_�����5�ng�������Zb:���0�5�8<\<��Dp��f��a;�s��h=hE�V�#��ҟL��� _@���%��9�-�����Ò�B*��|R����WB)2�EI�ޣ.�-���_�a�j�$@̩���	���e^�	k X�b%��n�+:��!l��k$pL�$��,Ҩ��kه���#����~����L�t�P�~T_��c���"'Q*�ҥd��{�J�TB��u��;�qx�!�r��c���W �F����Jyy/°-�{�ٗ��@M0'@3�%��F��{$��Կ���{�0�����^��F�p+�#�	�4Lc���2&H��6�'w�(a�°QO ��4gT'5��abd��`B6�n�Yt��:�y��,�=����J;*�)��Ƅ'���7�0σ���`X������0�:ܾy�W깮�7��I��c�?��#�
�&�6"q��	�|����������[�
�v�����U`X��]0��d��.$硯?�)
�3�0e��1�lޱ�ϟS0|���C�k0�&�4¯y��>~�G���r��/�?��g��?{t��w���=J��`B��G���p*�?�F༦�g��%�#?��[�
~o��O���.�D��إK��|t?Iq��7�w)���� ���;\v��A�^�t,6-�m�'x�0s\F�BKe,�+b1�9���(���u�������6N��jة��;�� ��-���Co6�E?K���P�N��$5�ޓ h���2����!*�/�\8��%���p#(XGD��yd�{z<���A��wz|3���9�ڐ��TՎ��Vx$���z�~��E�v)�7��ڢ�h�T��!pMi���R#,�'��-IҪ��U���[\l	�Iu�w�N�>�t�;y�O}�o��W�a����h�@VZ",�-�~�A�8��l��8���}�H�����7����'��:+W����q��w�w�m��\�xk��BEQ�c��e�.�,��	��'#>�	!	%�H*ƂU[q��K�?z3�Þ/>�����w?��w8]�n%J���!X�f���	���
�9UO-Ca�%$��8{�>��}��K��bGO�����K�p��y|��CL�`�̘���<�U6�ĩ+|�a��ňK�F���}�ڏp�����/�1f$V�_�[�n�Ɲ��y���xʇ�<nܺ�¢<�����^�;|M�$~�ň.�}�)DE�4\��g����5��ݸt��~s'y]ϟ��oN����0tX;"#c�F�����q��y44�ETb�	S�~ٰ d���P�T��7�����͙�7n�Ƀ_��ᓸv�~���}������u�/�:����c��`b�	K����o@�_#|S�g�X�p��n4���	���$��F<ĽaX��A	�-���e��p��9aϛ��3�*A��	~&�0+R0����|�F&$���0l&aj��<�"�fE��q^��W0� �JT),9/��4`������n�H*���Bv��u��ײK�#,���#��¹0�}3�9�\��;��`#��J���^�HVSu��4�cB��o0!W�[�=��a}�\���A����Q�����_�)�|^c[��)=o�S]�\%�&@k5�#�x�z�w���Ix�����=���HIT#�����/ 2�Ю<��ͪ��d�䖢Bf����)AA�d�0�o�Jm����״�S�\��~Ã��cR�%5ߓ�ѵT���:��K�H�q���(�zQu�Fp3�Bi�؈�(24�U�����z1#�#	�#��C�c�s�ӒρUt)�%��o2t�a�/�4Rh��J!�,��˰2X��ê`F(6!kaX_B!kR���j��r��V�����,�~���z���類�z��$0, �S���a�
�������pXI��NV0lUI�#w��@�2C`8�0�`�J�V���S�s�0��0L��J�� �Z	k�VA�����&��&߰6�A�(���a���5�z!�=`��f@6a8��$���`&���]�a�����~���=�<|L��b��|�|�d^�*��`��=��g�s��L5/@L0~I�}v�;��.]R�����蕩�e*Ү/�|U鹚j�4���L��N�o��T�]2�vb��|0�s��bʨbt6���1�Fc��&,�ہu����soZ7�0Ё��t�������~�}�yW�Z�%���M���*�[�=�`�w��k|k�1��J�Bp_ڹ��ɬGxI'B�;R<aecV1	!�Z>�����I(�HM@`�x�U
��+�"�r
B���?o8��/nv�f��7�`}���^A.��g&���|�e����$�}P�8�N@h�M�p>�D4^)���iU(k�/O\Ĺ�W�y���f\<w�N x�ǹo����s3S���'"�bq��=|q�,b�A:�C����?�7��/��'�0q�d�>}wn���Sgx���WG��gy�E8��L�'�?�ś1e�j��T����q���i\~���8+6�����詯���>��h6o݀��.Y� �Y�H��î]{����8��ID���;"�uI,@YS'�� ���Ėwb��q�1w&FM�is�`�̉�=�mM�)ȃ��J+j	�7p��s��<!�و�+E0�q΢����|����	�&c��7iazV�_�5�Vc񒅨�����%&O���?���{�#:މ�ʨRyf�;g����p��,]��m�>q:&���qc�b���ذa3���0�-[���\̛�ׯ���_�CM�H�_>|#��[��ԡ� L�&d ����S����P]\��k6c��i�:|<�m�At�vlڎ��20��ٸMC����X�l�%�;�����-G"۹�Tr"���l�XΧ���Y8���!�e�!�~��$�LV
���3��im	��#0,��%2"�yѠ���@�	d'�%U��u���Iq
#�HT�3��^���]p��	�"s���,C�aF�� �+op��#���Hm@`^;�i�
��FP�"cB�;R3>���Y΋�Id�����Y�z��y��am�4c��$�7$� ��,7�L�	��1�9�Hb�y\�vC��g\B�"�f�	�F���+�_��.���\�����TW�}�Ԁ��n����.�<��;#N�%\�P�����^bJ��,3:��;�J�R5�)�*H�H%��ن�3y��x�`G���j�;�)�>�g��.���<	�!#a]MC)}<z��v �8'+��YR��u���R��z��`0�D/��뚠878��p�{�P��X$��\�\�7�T��4HkaR��rN�`^�d|��a�9��;	Σ10h5�&�#xp��S ��d��E�:8��!��;�q��Jʃ+�['>�~�p�I��o<�*`G��'�He��E7��7�	���r=°�.���H�z������0�[�}��{��%0�J�%D*i��J@�@)��m�-�aK�����!�F|&���*0L��_���4���X���@�`�Y	����y�mTq���W��k�v�D.�ml�*��Z�@�aX[��A�0�b0�7���K���=�$��i��J���e�[��:���"�R�D]��7�^�_ �QZ�H@�`���wK��}����Ix���n.a8q�j����1s�l�ٸǿ����x�ϱ/=��/���K�ܕZM����ݩմ0��%�����?^>{�G�ύj��&$����2���??{@�%?缄Gh���k���	����Nh$�{�S����֕��{��g���=��`X�Y�k��8�r�o��%��|^�N��j�pV#fN�Ęa9ݖ�ic˱pf���T0�c�l|�c!6���YӇ��,���x���0��>��1���3�	:���k�w-���w�d�'�����ip��أ26�\�&Ws�N�5pIi�k���RiC���y���:���g�xg��o�h��2���J��/�6�p���#��,�\���Q	�@v��Ĭ�i9�e���}G@�h��S
(�"���O�o�hj�d�cQTӁC�/���K�7w6�͘�mmŧ����C�{�;ܸr3�L���'���?����o�ı���U;�$X���+4�>�? ���q�WVbȐ��2y*f͘�y��b��yظb=��^���<$ǥc�ރ�r�	&�[	���F� $�T����a�������Whَږ:L�6������f�
:t ��ۍ��
$'&`Ϯ�x��%>���2`�	��,�yE !��	��>��9��쏌��V����m#Z�h�|�{'V�]���:L�<�y���Ő������+>Ai��d3n?~A��
+�PZS��cG����MX�d��ۋ���"&&��y&��l�u V��4v��A@q�FA�8\����^@�СFBt"*K*�|�R|��C���[�$(�/+����y����GEu|����B�WL|��7t�E\A.ݹ��wnc҄I�Ä�1h.�GIz�/Y��^���'X�x%|�P�_�˗�����f.��{�=c�^��r�Q�%[��O&L��aB�q�*C$�x$\c*T����q�l�A��|� 2g~�Ҡ�e���K9�p�y�4ye�+�A9�*�G<���>é-*fT��2�J<������@lVD��V�i����K�0%1�\�gX�mt)����Z�{�t$�3�����.�}�x�*,��dZJ8����V�=�a�V�j0�H�,4���=���J ߌ�$��=e�O��T�iD06�u�) �� ̈�CvRo�e���N�_}n�O�T�����Wl�C��	וL�z^r�s#ª�!�\n(� �O�����~~��k�A	��a]��>��l�F��۫aפF;�W��F<���zt=2x�������h�,�����OG���(s8t��t'���W��|��pY#>;&��0���,Z*�U�&�
�<7��*��=�C'���ʶю>��0��葰���Q���O� �c拿8����o�¿��;&�x��
��l��=#{�3�A�A4D��ֻ&xo�3t\Ra;��>�g0,�S �
��W���{�����0�[�}�����O#4S�2��6�D�e���~l/bL��h��Jܴ';����� �	�"1�][D׼Á�n�x��6�(N�he{1��~áC����z���~�y�����HA�&��/!W�J�Z�q^�a�k��_ 8��K��`8��#3yM�UT���zL�6��?�~p� |g	��a���amэ?��?��w������޽�G���!����xB�}ʩH�0a���+H5�gw���S�%���e � �&t�����x��,YG���F�H�Q���`����
�7���ՋGbѬ&|0�f�z�`��:LY��#
1kb���e�:�j�hl\5;6@��)�QV�G;��λ�_� l�},���qC_#O�k��-���: �n�0�M��
;�T�X��R8��/����D���
��v��6w8�
� �p<��s��J ���<�p.�8�>��e��W@P&L�rB�a��-�\��:�3��=;+B�87·��V��+��ţ�c��
��G�GQ�7t3��sÝ8v���:�B\dt8��0n����m���q��aii���	���F�;s)y�~�T8x%�/"�=�������CC���ƆFL�2ƌǆ�kq��1\;sS�LG!���c�r�&�Y+�T�s(,0n�\�u}�YE�HHO����f�*|�����8�>}��/�`ӆ����T0����8t�4Bb�a�ٯ��'b3
p����6q�T�y����
��ǜ���x�B�����}���3466a�	8u���>���Z�@��v.�1w��}�O��I�((/�5��Κ��������x��!��p��Idd�c��x��?�mߗе�BK����}� dV'?���c⤉H�K@eq5���7���x��1���G�޽�e�
���{��'���ja=��p`۰��K�����	)��t������c�����0	�,Ǵѓ�g�n���G<�V�؈Аh�����%��'́�G"s�]9�c�Q=�}�	��	��mCx�0�Le��7�~*B��	�y�C_�?߳��o&����S���0���Kt4"
Fr��́Oj+��F�6�pDȱ"pz��8D��HB�0�T��Z� ��'�������Tl1��kS��_�P��,���7J,��Z�<$��)�ǋ�QP��ώ�<�.�kr=ܒ�N��:����Q�I��ͯ�#�E�=�Jk�Kr�b��Ih�3�&�R�U�s�g$�&��D�N�)�$Q��c"������,�U+�ލ� U�_�n��<W��}r���Ro��V�9�9s�}�)�gXR�"����!^g��^w�V��aj��|�D� ,0,^a�:��" o8|��I�#HV�$��R ���f�\G�i�u�P��@��e�B�v�� �|hXZ���J���w��%����x���a���ѰL���:y~��g� S�T5O����1e�
��� ��/��U�0w�:�X�ӗ,���`��=�`�,X����BRn��,���T�S���ׅ�p�`��w��������Do�a��&��+�[N����{NI��L��v�
��sIR0܇��n�����A��3��]�{�&�-k�&z�FO9�����j?����=�pu`���_��wiP��? 0�0\��<D�����n���W��t� |�\�UֆHk
�i��g���s�:��ܾ�Ҧ=�w�0|O�O�P�°a�����o��)ɼ,��@�&�9��T�o�a�U�F���5�=���4��a��&�_����0gr-�Oo�6����w�gb���:�dF��h ����O��_o�ﻃ1��	a�zz.`��M�����,�`��H��G��7��	1J��NegOhP�V�R�J`Ց�K;��&x$6�[�͎އ��L���������$�g��e�4�raH�U�/}[v���p-�kH�����V�i
/�ET1,�K�2XF��J��E$yX%���/�V��L.&d~�#'N���^~^�+�#�v`��i8p`~��)����^���`h�P|Ƕw��Yħ�*/�-���l��^����.n������M��d�"̘2�|��wؘo<V0��Q�ݻ���`�ܕ�p����H��C��|1n�|\��_;�Қ
�D�������đc_�ރ���O/�������E��CH|B���$eU��/�!)0��FQmNw���W/���'*�*��WY$�t����Gq��]�nB��U8�
n��6z$��|ad��8|�x3�<~��ǾFJNR���0d򊋑�����/��������������������cе��;R��7}��W7�^���@-_ j�ia���%��W������7nbŊU���eǹ����n���m�3v�ɰ�Ʉ�K*����;5��������s��ٰ��E{�,�`�Rr�Z��gdV.[������rFFz>�=�kW�a����GN�0�w���=��}���h��"""�	�U��B;>/>��"�'X����,2�%�6�i�&L뱳1��V�a�ag�v���#�`T7[��+�IoS^J��_ �8P�U�!�ZE�s�@�[󜤒��&蚉�K��] ���|��e,�a�D� 5	��_�#T�.��rB`![���20�6���P�Q��6F�U�&J�)���y�9I��'^_㐟{�5e�%~�X�g!�f�U��f^�14!|����rm��l�uy�WX$�]�$�AB+�dJ�Y�Er���7����g	���ӧ1�Op��υ�_6t�l�Ozg*b{,`'���OW(�@�V?��}� (�A<σ���G�w@.�8���{\O�}�AX�B(�P4
��հ��d�\C�K#±E��Jn��ha����_&޳�¿���φ.4؜�'}'���#���=��`[�Y�o8�=#g�����uŻ�x�:=��S]�(PWOm
�a������g/�臿��?��|��_��;Ϟ�՞P_O��Wo?Ŗ݇��8��H���`X��/0�5�K�D)�p�W��	�o�]�C��`�H��	��w�	�]0,�a	�P���f^�[�2V�a)d���0�0,y�%�����%߽ROn"�t	�J_-�W�u
d�HЍj���6����������į��+ ~ÒM���>�C.A\Y#������a�g{p�ֵ^a°��W`���/�0��<�sO�\�����:�>���~#,!��Lexx��_<�@�������]/��]-�JXD���7VX�_��C��ź�0oF3F�Ƹ�̙R�U�b��6�^Ԯ���)��7�g��y�X�h4�-����PU���_�p���������}`�@#��Z��1@��0��6�0���w����hNX�pƻF6`�3�`�r8��B��]��;Er���#B�	"3v
�$,�YX��a��؆��M`��Y;).�@�2�_J�fÎ�;gv:.�pܹ�!�>H�;�pC?I4�@�5:���qu���J:����k?$�����s8s�:Z��%���@#as���ػ�#\�tgϜ���3��′�ܼw_;��DB��7��"��������q��1$'' 7'��?�<�%E�3|���8��)��w����pww��Vl�s�@\J��{L������}T�.�u�GD\8�,�Ǎĥ���O/p��hmmDjJ2�}-����ѳ�΂�C�*m����\�u���+7����+�3SP�L�����?w�ظu�*��菆�F��Eܸs���04�T���,܄�O~��oN #?��KI���W@���a���7o.�b��;>���?��8�0��vA�0�˳�m*�W<w�j��ao�`�0�%�#)6��4�--h61����������\�r5ͣaCc��3���0'p��fb��R*�p��]<��{̙3zuacb	7�����&6�0����e�
���<<x�e�G�y�H�m�gX�0�yO��Q��H� ��7��7}m����-,�C�n(�Jn@@�Pĕ��_;/�MC�x���#�0��.�W��1vτ��I_6fU���<�W�0	�V�P�Q	�x��A#)o,SI?� ��X�œl���畿�%v�&�BړP�(�.�W�L�%��%�A�8N)Ӑ�
&���5Ҝ�q �i1jy,�$��Y� 6�'���֭A4D�}���0s��L-lr*q��ya� $�u)�F�xQe�xV5�~.d��|�O��)Mf�.���A<OJ���h B�����瑆>nRI���Cɺ��p&�t�}B�,�!�
芧N�[���9��/E4޲�P����63l&y_�i���يƑuA8�zQ%. ��0b;2	��]Xۥ@�.~q�H)�Gi�(T��E�q�霠T�:�um�6��\?tJ�G!���[N+�&L�a\�v���6����EÈ98���=q��%|�o�|��7�W��d!�o݌��.�������=v�Ju��E��8oKY��J��2�����.���o�����O��7���N�{���������GX7������/��+A�]b��ayF�T6�w��W�X5�N�i�=aX�Al�b���PT�a°QL�	��%�3����o�G򹈧�*�_��!�' ��w	��᠞� q7˿�W���0~�k3�«0	�7��#�	���Oï{����%���+"���.�)EF}'f/����b���q���W |E�]�e°�c��`��s��=<�}��)"��%�
�>�°����r�&��H�%k�
�{���8=a�)�[����c��&�hMè��1���`͒�_6���ܩu�;��0�J� �¢���0�u���L��Y_���*װ���020�)����ka�+W��a����}�����j$d��/*	v^܇�/!5΁�p��[X�BS�ip
J�#A�!P���K�p�Q��-G~�Ć���� [������s`Aص��e�Nԉr����JHv纮aǰ�س	�0N�YP���e@�`�k��՚���O,<�`��x�������[h5
VNv0�6���.�SSCx�� &&�nx�������^¾/"6� �g�h�'b׾x��	.�cb"`bd���DDGF���a���/EJd2,l��#G����`᚝��J��{(�|�a���	���q���8v���a��И0G!2.C�Ų5�0c�T��bc�q��1<}F@%��dB��>1Y0p�FB^.޻���;�mZkµ��#����3[S�x:����֦*g�aCU��k�nb��1pt���U x��������G�(�rt���<��a��N�������4��ضm'�`ϗ���+Fn�p�A� dT���{�p��Z�����۞�)ۤ�	L��a)%��m1@g̬�0냹�}�)�]����l���K�(�	�UE�����h�2���c������V��060àA��_F|\\}��؆'�����X�z;�����
s���Ap;0Bs� ��M��1���d��$�q���B��y$��#����I=޵� �X
�<'@��a��ZD��Mx9t�3�v��x4�١ibU�U��Hbj-�7�\��&/�U��=@X�pP���(��t�y�E>��T+	�$6��
��ء�_��>G��r��8�)��)���[}>��"=��Y������$����MZ�}����3T*2F��8	'�8a��9M�/��ңdЛ�xj�`Z멕P��I-���s{m����>Ͽ��x�z�j�]��C��%�ܟ�����ɶ���gZ�
�x�V(ѨW�:O��@��%�x��w���Z��;�m���&Ex���v�еMA�0�g6b�G�����xB���%n�����<��ox��{<|�O�����������C��q�R���YX]���|��y��c�"���G�9�����C]�9�!;?�M�(�(ALJ
|c�Ί���q��e�xU�f�"�BU�3� ����k@�g��ޠ�& �ޠ����1z�j��D����}������� :4�G�3 p�5c�w�rL�;4�$��_�¡�0[�a,�6�	K�a�k=ĚtZ�H��L�u-�6��0ܟF��c	Ñ]0�;ax�����s��^��`X�į�0a� �-�)�Ѥ<�*~X<ͼF�	�9k<�?�a��;�s.�@>��I�C0j�xL�9U�����_��˗(�gX��a���<�G�s��y��I`$?'�>$0���Y��kzx��>��_m	�w50� X}����o��A�����֘���DL���s�q�lY=kw`��F�S��[�d~;�/��3�`��b�4f�0/v6��������_8�=�z��000����0HW*��<���"��"&9���E@dB�R�O@�
��gH�������Lx�e�#$��R��T�+e�#0[��r#�I���Bv���ȃ]h.샳�D�u!�
��ep>��֞��%��G���nT>"��$�`�
��B�+��1 �nHȯ�G_�����a��p�� Z��њ��)�����@�<�:�@G [�p�����#(,k�˽>���|��~<z������!x�ݷ;���X_F:zp������	éI�8��9�|,ۼap�1��+�p�j8f,\���8��T65���~������5,��7��"	�_;�����ߜGrn�<��H@s�@dN�\�����?�	�@oX+�"`{�r��v����=||0~���p��}�i�f"$<	����~a�?s��p�����?�b��	ߠ��!.!���HKM���?���Ga�����8١;F��y"�>�.ܽ�)sg":.!~�T8�����O_����B����5�6���g8{�.��`ؼ�wpEa���;xH���a̜9�'NƤ�1}�L̞=-ǒ��r�V�ߴ�����q��-̡a"����Ca�'�g� �ވ��I�'��  ���#�������=³�	KqB�a��m4a8N�E*�y3�gx�{:a���3,0�G8�°@�x�5Y4p�:�L�oK�|ikaXm��m�@��������zf��
���2#?��x�ՠ�.�m2�L�E�T�¸Q��!�.��7��	��9�hwI�e&g��9I�&�$,�)�^�0K��
�k�%�9Q�&�G���R �Ӽ��, �@��1��V���'X�j�JMҪ��LS�a��S�J}:����)����C�q~��^���Q"��#,��|��	β�6��AXJ4�!��u�h��땊�\��(>�0r�P�d6�&�����'N^T�+�|��l�J��z�Zlغ	[wl����p������ø}�
}�����8�f�&�n����Ъ2 ��Dc������c|y�ҳ3aek�����d|}�0nݻAH8�ūW�+"
��꠴��0|�=|�֙K`�w�.1�8Bo,�W��/z��0,P�4_�7 pO�\���u��-�޾��o��ߒ��(M%:��f>Oܟ#�s)�ڥ*~� ���;&V
�D�0��_��b��tZ�:$DB�ٖe*mM��GU�Hi�1aX<�o�a��_��Wa�uIH���X%w�ۼ
��y�.�.�&�
�Sk������	��y��50�&�U��w6�߄��iaX@X�T�Q��@eJ��-�ؠbq{�e���=%!?aò/99��	AX*�=���0�3�:���7����p�����[q�&fX�$���֐@�a��,,�]�mk���M��i�h,�ۊ�sg6a����Q�=��ۋ0�5��qp���{���4�/����?���>}���E�1x�>LL-	��ptu�7�$42
ށA�0BO��	�i�����?�	^�~Q�8��q>n~�p��2�T@"�K����c	ah�{q}��e��h�],�]d�8�/[vb��,��EN�a��tX�Æ�mC�-�c\1c��]�"�D\�U�0����	g��غ�8���K7�@�Q��M�?u"F��1�a���9a��[��}x��3?CGN# ��OH|BS��g����g���6��\�q�aΜ9X�`�/[����=X�%Vb���زu���מ �wD\q�R�����X��cҼ���8w�!��MDTZ*Bc���P$�!��qi	�+�'���9A(�G�����Q���B���7q���I����S��q	K6����0c�L�ڼ�Z��[Vaۮm���,_��}uX���|�3��Btj�Q.��*0�.�y��߻���}��+7`���ظ}�݈-;?§�����رcػ�S<x�w������{t��y�������ɸ��q�G�̵[ؾ� v�=�����C�q@t�k���v����]�߳S>u�*Z���=�^����cE��20��	�U8u�/������x����o�������ç?�����i��;h��ę[2|��#a��t��r�
;����<�g����r�"�0�[����x�,��9�Jl�U�e=v4�95�#�L�r�i`��@.w��EX�(��
�,���T�nɏ�-����@�����*0,����P��J���$��9�gX�*��*�T`Y@X��R�M`P ̘�+a�	6@�V,a�`��6!���aY�\�R �}�#=���^a(�(ka؈ۛ���m�+�ن���J6Q����r��
(e ���L!�x^B����z��Z����n�N����q��>�5PL V ���e�s=�M9~��J<w-�ˠ=�}o�Ĩ�x�=h���/'	���"v�����@��� ��~�x�#�8Ū"��^��EB�,%U��[�oa��HM��	�^���A��H�e"/3���>m.]�IcX��x��}"0�����~�5���i�p��8z�[�GG���'N�{�$nܾ��O�����s�sV����7
J��剣8~�
�.�QT!A��C�]�!�I�f�IB;,SF�4���#JP0�.��~{�7���ס�g�Su�7}ߥ����}o�U"�#�v��u�KLlt(��z��tjؾ���c.޲�}g[x�m�3̩qx��kU%@a)#e���R�h���ۯ�NH�ԥ�h��a	���|����0	-�k`8�J�ۖ<���B[�)ֆJHܰVo�a9�V��*�@.A���\ X��a��'���	��z��  ��IDAT�%L�iu�&E7��R�����۸�� :������=����:5����3,� R-��]@����������@��� �-%Y�`� ���e��0��y���&-����8yl/6�� _}������۱m�̞\�q���hN��!��5���O���p���عi*�L���E�;{֮����:��V���d����b �z�������V�04o���=��� s������m�CQR^��`88;����N�
�O�?\���UT��!C�;w?�Ĥ���w�x���ɾ1��8x�E�����~p�r���|�}`Ɏ5���T��#@|#��U
Gv�Δ�U8�#�ɁV#��3�ֱ�J6�a;°=��1�P�t�·KT����T�u��c��]���'ù[4>�?ƍG�p��<��%�}�w^<�헏p�z��c߱o1t�<�U�CR~|���~�;?nji��<|��?��=�#��\x��\�n=�n� ���~�r�̇j;�r'�7����GL_�3���g����q��y|x�sl�t>>��:�-��=��N��qNo>x�K7n�Њ����}"��J_��k����l>|wyn�^>���9Q�������{x������!�������[�ו�?��[�1n�DK��N��4c�U�x�	�?�k����=�������%���7��ۏ���!ȔxJ��.a����d�n�Gg�ʅAY�0�MGJ�h|�����k�k�]���k���=�1��u{�������g���%n>�n=�;>��J�G�8��gl63��Q��J؆�!��S�o�'���'8}�*�}s�p�O��1N�������/����'q��E:ym���3�:���Ɂ;��D�1�!���p����
�	����I�JcE�qO��s;#�T���u&�)�, lF�!���@��}f�=�A��h⅔,�IB���_��FL�X��ځ^=x�T��EW�P�R�����%|B�XB(4��a�"K�Bd�
v	��6�'��MŲ\$�Tq˯��L�}��D]�_�Bd0A������a	70���3,0,�"��"Jǩk��݃�$��	����$B������Yoi��mĨ�B�[�W*�2%�UQ��H�����u�^q���r��ܗ>�^�g�N+CJ��H�H�\�xϝ$��OBa��a"�\�A�X>+�%�S�EO�	�`�'���ї�YB�@�d�%\;D��y�3�J8�0q,-M���ٳ�a�X�t!vnY���������:������gq�1��m{��R
��r�&��=�va<?�8�8���se�&��a܄�ػ�S|�g����/_����8q�<�-^��"�6���S��͕�(꜊�<��2ĵ*�Ƕb!p ��X<�%3�V8�i�!U�������	���T��5 �	���`U��&�U�?���{��ð�%_�І.�Su$����ҡt�j�Ϸo9$���qx�9��X�� 6@ɿ�����sm��Sy��=��-EUD|�)N��b0��|Oi�)(�L]9�%tb�;R1�"�	1��*���@��^3<�=��W��0��B�E�Z���@�
�Z� ��g�z��H�W�%Ӟ�ْk���$�0��EL1a�S�������~�f�:V���kz��l�����9a�a��@S��Щ@��aX�h	���/�p�}h��a��	��	�o]R@,!������`��r��n&q���r�sس
g�cxk6*��T�a�*�ں�#q�ӥ8��vڷ�g���"�Y���+PY���� ��x���&�}al�~~��hoĒ%s�j�R̟?|0S�M�\���[6�T^̟����{�")=>��H�NU��,���W�{���>~
�,Y�-�|��{�Ħ�a�=شm?6n݇5wc_��6�@����-���qmX�y9��ُ��kB��tm^�5�͇%_�NR,  ��¤l�cT	b*�"�y*�'#�b$B*F!�Ӱ��(�����4��EC�T���j�\������;?��;�<_��=��\y�7�������̝8}�>����x��}����Ȩ����N��Va����:�>x���⽧�t��E��2��{/b�F�ܭ�8q�����Y[Y2~��=	�I����AØ�}�6���;�#^!D^��E�޸����Q������ܵ��7!���q�����3(:�C�P7��B�1n�N���o���[wp��#\�}g�_ƙ�.����؅K8q�N_}�����G<�ik�"�f,|R[��ܦ���g��o��-۱|�G�����Wg	�O������<rG�����`�1s�*TwNF`j)A���'����mEՈ�蘶���b��;3&-ڂ)K6c��M*�Ҭ�0e������~�LdUu"(�>���5�!H�4"(�NQ�l?�j-�)ՈK�DV~2s������JdW"�J/�@b~1B���p�ֱ0�I��cl}��܄���*�H��4�x%�2�ӂ���pK�U%�E��L��s`N�1%����%�Mx�R����0l���`80��Q�璤�ObG=(�o�XU�+��}�k0�w��I�>tqd�� �WX3�N;-P�'hm�7Xk<������u*	�ݢkH)���p/	 �w�3�B%h0�$�VB#�wK�lh�h?�W�h��	w�=qJ�W`lO`v��_\Ǿ��~Y�uj�� �V�"~'�{��;YG��n/#�m)��������d�V�\G+�.IF�a��, �^M8�
ϠT'?��� �8w�?.Q_L/N	4��HXEt�������8}�".\�����!77��ũ��q��ܿs?�x���C,�;ΎvHMM���q��߰x�^x���*�B�����4R<��<n&������Fyu5�;;0w�<B�D,_��}�:�-����S���&9u���E�
]�)�p@��-�X)�
�ء0O�U�HN���yza�fw	g�k��M ,��=%ߟ{h��2��_��i_=�{�7�0AX��$���j)��VC ��j�5<�Wz��WG	���ߚ�j�J9�c��=�����D����ERQ����2h� ��k ۍH�cL`8AÃyo��}�k0<(��T�/�p��<���X��=�2�����r���pO�q_������𶤭S0���TD�&i`x���_�T�;u��\8�@��°6��k0��� �œ{��X��G�W�{������[��@��ðx���ab�*�0��3��EZ���-��cl۴ ߞ؍�wN��z�x̝ڌy��pf3�N���q��:���jL[���K�R����0�f!-���6p�Ӄ��.�m�aa�[[#z`ذFlٺ_܇�[7b��5X�l!f͞�)S'b֜�>�#�G[G��T������T��w�����]� Ú�[	�{p��c\��H�����|�)���Ay��|�K7���OIcF�����K8D�x;�����F8K�4�LX�d���d�pb��P���Q�o���!�Q7>ŝ�-�Q;� �sR4a����J9b+;Q:rʨ�Ι(6�3Q�>u\�<~!�F}���Q9jʩ��	���< ~YR5o6��b���n_8|:*F�R�����i�;�cf��}2j��Ω�>�m�]�s�o�O��'N@@�H�%Er�$4O\���b溏�h˧��n���W|�鋶aњ=X�zf/ކI�E�vcܬ�霏ȼN�g��?waX*B�z�D|�ėCj��w"��YE�T���DH�ϪCBv+"R��1!Y4Lԑ�c�7���1��O$<C`����L�T��S��
Wooػ:���F&�0�����������8
	���<	=�|�څ�#o��@��>v��m�{���z�}���Q �B1�8}��?ZE��/jk¦�OL��a�#/~�'�y塯Y��ཁ���1�-|�o�]{���l0��
̭�o�={g��u�]3�R��ԡH*�������5^y��"��T���N���B�;z�i�2�RZ�6��,	�R�y�st]	��&�����9�# �]�9HG%U�40̎�5��f.!a������a( .S0�P��J����b���L��^O�a�i�c�,6T���b��EѪJܯ)��g���V�]�̘�k0�߭<�<���5��
� a�( ,��dp�Ud��{֊�����x�d���F����D�$��J�X��ߛ$��:*��լK�b�H�sx	a��%����Jm��.)�$lB�)�ʚ8fM�aY.`"��Ļ�'׊�^��Z�mN��.�����惻>��q��<�ok�T��O]=�K7�`�H�HEAA.&M��M����p��aܿ��Yп�����7gU��E�?%���P�4����Fb�c�:'���;�d��(��@{G;6n؀�������q�����9v��R`���r�<��~E|��<0��P���FzR
�F�|�da�w���H���ڒ�m�y��¢ޠ�S��ߴ���0J V���Մ�*~W�����s
�qJ�{.)�+A�/�DX3�)0l��h �mJ�w��c�>�c}�z��x�%\BJ1k`X�~ls���1
��0\�*��ς��%a��}0�SZ ����p%a��0�K��}*$g�}R��z���y�>�lؾ�^8�<§Ξ�Y���.�����_õ�q����7z�k0�\*ωgX<�
�	�XUM�T�I/��X#°�5���g0��Z�7X#K�u5pN�%vX�ϩc�����_<���wb���8}b�^?�/�o��US�|�H,�=�O��US�j�h�pF�в�HByA4
2Ð����� *����q����-��,`cmD#>>#F�a��%X�z9>�x;>ݷ���g�^��k>��v���6�P˪�QX^����h֊ʦz��cΒ����#���	��ۆcg��}_c�'_�̕�ض���߅�����7g0e�|�ٹ_�=�IK�#�r$\�J�)!Rܣ.�e0�j薤Rf9�rK��sr=�w8�+���t$<�����k�w�P�����,l�_�8$��%��5pOfgEx�PD��"�F��#��q\'�n�����WM@��i-^����Ι���i��i%��#0�� _�}e�s�]���
xDf�-$�ip	K�Cx&l"��N�	(�����$���BP�p���x.Ep��F@
�)"��GX.|yξ��ʀ_x.��H�OD����#Q4A�Z6Q5s�����$5 0��)U�/Ddb��K�4����&>��b��܆���ʐ/��v�,��.
�^p���?����Z�S\�N���6p��@tb�bc���cK�Y:�Zd���:� B#��^����h}�a�{���LX�$��9v|�ۻ�{�4ػe��3v93v���y�G>L�	U��aQ!?��r�-���g	'�8����?
��ap��%��t��kH��;%ǰpφwt=�
� ��mpA6S�h5Ʌ�В���n!�` ;�l�c�C�Ҵ!�`�E|RZxNY��o��%6���!j�$4�a)K.�}���V�ϹS��@�H���c%	�
���x!�*��j�����_�y��7���4�`Xr�ʺ���R�P(�>̈́@l��.�b��.�a	qx����^_fD6��ྻ�^�^L�%d����0	� �T�zHb$u�;{K}�ɾ����Jxk�+�T��7H���c��)���+���m��#�3&l�o��%�h�/�2T��$D�S �:�Zy�-�4y��D^Q2��(�V�u��}|=����m<�y�t���8{�-]���*TT�aԨX�bv}���݅5+�"���ӿ#!9��kO�������+�md\���n[`�����q��O8|��i��iSp��8��1�8�%�}y�6��w��	I�����|v�(����!�h�+	���R_�2����2\K8�֡�@�I�0w��/��`�p� q5UI8+C��햮��}q?�4Udc�����6�`��/�7"	��,�8�+ ~3k<���"���?۹Q8�	
���ՆIt�V���0�@X$��S�i=�o֫	��W�K��x�b5S%���)��CjYOO��j^�C�nOϰ�p^�g�u��`>ax.ax+N��Xש3gp��y��߂� ~��	a������IP�����
�ˣ�[
p_���]R`,�
���: �Y7	�Ěk*���� ��S%����Oo�ȡU��ѯv��j��~D��)cj1zh1�����i�0j;&�Ťu�Z���4gǠ$'%�	�8BqbC}��og��8���	��A~A&L�U��a���X�j)6l\�m�7a�G۰㣭شuV�_��+�}�P4��c��5q�뫑�����d��c��h��I,���a�ڝ�0�W}����[ف�?��K�q��y|q�V�ݍ�N�h)h]���8E ����R�5�N�%���=; ��a�+��8o<(��6%/�{��'��3{��Z�ͩ��R~\7��	��P
�i'��3�/�`��u��y����L�ۘ�*\���y��J��O��k5�)��b�f� �0�W���b��j�2�V��{H�Xxf��G�HdO@@�hn3�0;� ݎ��zh��
�idf��]����L�FtZ5b�kH�!4�IE�/��/c8<�G�-}�	�n�	X��;��+��0\�8�7!��U�X�v7FM^���	(k�����"̕�#�`��fX�%��/YBR�����\��Z��}a����ñs�.|y��}�:c6�+��o��R�BV41��p�)�Kd|h|�#b��k]���z���!<���9AU�c'��_��8C��p-�Ch9�c���ξ�FL+<�Ҡ�k�ψ��hP�8}���Ϡ(��O�{h$�C����r^�^����#�r��\R	ۙp��D�Mt�xg6B	pycI�	��@z�,��9����Q	��rJ��oL�3V8��i0"d{�
�i`�Y��^�p
;a1��P`؟0�O# @�����f�'�K-@IL����b+vVê��XSX�'(�/Y��z�|�+�,���L�;m���W^a-���~���C	� ���h�њǜJ���C웣���`8)x�[E����� +��H.���h�H X`�[#�����$��K0,�,)TV
ٿ��3,iԴ�7�^˵�&;I%;��I�0����x��ܘ�W��2K��i�d�|/�l#h���@�KAvM3�9���ż�1s�L|��S\�z���=ܽsW.�ù��`��N�#(4�;����E���!2|�\��)v�a[�F��p������q���c��q��n|�ŧ8�{'>ݾ+��@s}#�*Z���<�ؽ��>���3ض�`B���>�G
��qT�;�GB�^xLb���0%�D�) ֆK( }�z�jO�_	�u������5��k#0���[N����4�qL��6���>���H�����%��[2�sNTq�&���ao�a���a�WM㤘0�@�&Gq��_��>
�[	ÚX��=�?�@�t���_b�d}�v�����~_����l�z�M���c�{�pC�,\���;���ŋ8{�a�,Ο�@��`���a- k%�n����W0,�Ô������n�7��d�x5�u����?���c�?��M������w�q���X:o4��e��:mu9h��C[mZ+�1�6�e�(�MBI!8=9)��HERd ����� Og[x{8���@X�bc�����۰x�|�Z/�u��f�Jlܼ[	��?܌I�ƣ��
�M�7e��Ý�����h������ђ~-,�f��71c�Z��ס��)-���CI�X���n|��q͓� ���Y��D��7���&�H�ˇӌ��U@>�C��ъ@)�\:�Y��v���(& {�2~V"`xd�ɔO�0�J�h���-�q�� LP����6j|�	��	�s	��7m*2G#�`����q7wo�u�'�/&Q%��x=f.ـ!�g#*�
A��-"�f�ʥD�d����"�0�C���z�W��t��wb�u:a��Faȸ0k�f���s5m>a\7��q%#��玡0.#`�8�/�D�Fa�l��LE͐�h���1u�R>u����������0f9ϩ��YOcT=�	]�AR�$v��ȯǲ5�1��o���|��!�{��_�çOq���i"�����)lA\�dchDL�p���(�}J�A|n+Ⲛ���R˶�%v����U����,�j-�g�xς�xz|)�����?�/�A��|�e#9��%�H�(Dza9�G����k0y��r��xEf"!�FI
�Kd�Kh���;�0[�6���@�3/v0�Q��L�6��H�*�~\��aA�t���e`���.�]�,B��$�3,0��v*q�}�aɀ7a),��c(����2�.����D�D$�@���U*�@�K��xb)�\��4����j�!0�#L��X��2p�L����$��0����_�a/�5 ��a���F20M�9x�Bkc�E�tj����xp%�Z�E*��xz_S6S�ht�TU�뒬��Vm/1��S:�`n�J��o�@j@��A�]��Je����{��� vJ���wZ��,!%��7RE���h�
x%��s{#_^w�� �`dV7���oq��5,_��Ǎ��5�p���8��A�۷;�o����0f�p88����}v���ywѐ͇%ۈmt=�W����Ģq�t\}�'ϝFMq&&��ƅӰ�ںd&V���#�P�����l�8x"!1�|�%N^�����	���N�l+�aɘ@���=O��l��@b(��q����������E��������k{��D!		�[9�s�B(�A�s6�q���M4L�9pXa��7�[4���Z{�Ͻ��U�]]]]����ɬ9;X�j��M%'�Ü�@p&�>��U�VSbט��)�ǯ�n�ϖ���_� y�.��_�a��1-0�nf��F~fL������+�k�y�W�,��z?�؈1.a�w(��aS#>~�����a�aս1�I'��З ~�/o��-��S���`8�N�6ñ�bx����ǰD�<�?���0�Ga�21|��%\�r7��kz߹���j�1,�%���ϟ����'�LBp*p��0����7?ʔp��1��տWp+����'z�o��噃طk5.�=��7��ԧ;�s��Y<����I-��Q��ë1�}:�j�XU@��P����dƇ"/%�ɱH�C���<���@���S��Ҁy�fa��EX�zO��{�v�p?�o߄m̎�[����X�v�O���FՖx�¹�܀�<$�g 0,
EC���Q�f����X�qqS���
$��#0&�<�����<�{>;��a�H(�%���ל�
xa/B`n��;ߊH��TF�s
-�Kd��+�~"�L�/�+ �#n���tq<��k�Ë�o�+K$�A �	&��!DpH�݆��D�� ����͈�|Q�?9S�;����i�HkG@L	���p��m<�#�f�~m�:QQ߂�;���ۏq������y�"�ͅ�/�����|<����Hb8�����(W�i�<�;�9�>���?�ɫ7q���O��޷/��/��ŗ(k���a�g�C(�/�W�H��:%բl�|x�!.>��<Žg����g���*��_����^�����s�!��p���h����E��7,������U8r�ߵ�w�í���я�������p�n�GU�Xi��X
�J8���A����C���.�gX&<�R��7�N����xع��;C[�cD�,�'��qp�͂3c���4�.���σ}�G�d�5a�:ן���c��}߇8r��=z�G����/6�� �Ee�k���B�����#��\�����^@f�*�#X�(��{�{%��/Ҷ=��9����IܮJ����x�t���8;`Ƌ�!�Ű�<�g�nѤf�1L��U��MXd�D�k�x�B$7�	��$�7	�w؇����D�.�$����Y��.���{4�Tڙ
�et95��Ӈ���u�o�2�,�}�9}3	i7��X�aX�F�á��.�ʼzL�6�D���h��j԰˿c�W1,�Ԇ�s�����8T��Z<N	u�I��&K5��w�DA����H�ƒg�S����b{���m���ɫgq��m�Y�Aa���G0�Q����EXH��PVT///�F��g�q���{g��@��Vx�̓��D"��������;P[�����X�Y��#��xl=&+@Gu2����~FVpu��䙋�vۇ(l��h�Q�� D�c�a��A��9�bI4&(��Ò�$��ݰBpAK�J�D�V��-|΄8�)����6���D�Lu(�'�$	īD�en�)��)���u�:d}���g�w@�m�s��O�!�{�Uᵀ"����#��7����`��\�`���J`���1���x,�E�t��>j*�dg��a��[���1,�$�fX0���Jbذ7��gb�"!|��\�x׮\�͛��oܾ�j�o�w����=cX_3܅��b���İ���aX��=��F�G�U��faK�o��hk|�3~!���=����c\>�[�0|��	���]|������N�<_|��nű��޶�X�t
�Nn���r��@uQ"�����`�G� >�����
FT@ �BC�:lV�X�];�����kV`�ڕX�^j��b��UX��Ｓ۶mM�1���؉���?�'�~�-����Ή(.����)H�( '����X�a�K�R���V��ף����7�����70m�j���!�hbK�V��
�5�;��H��?h'�<	a�aH2)�f#�vK��:x�_>�W�Iw�&0������1/Kt��v?'8����Ђ·AY�H����q�+-���˝����)��ȼ�ܞ"l��	�|�>:r�>;����oj��z(Jj�����x�#�d�~�d��?��S���-����)͟�pb8�h�|Z��;���)��� G/_�E�p����Y�x�m����^��7o���=k��+�/�	����-��+SǄ$TO��'p�����/��o����5�8o�y���&����A����Ϩ��~	��²Hd�ɿ�&Y�C���8}�.�x_\��3�/bĸ�)���;V�}Wo?B�%�����wz�b�g����20�9��sf���
IFPT�����ÂU"2��Қa���!9�%��a��4��'�"0��L��J�3`�+�x��y��x��ܞ{x���� p���߹�:��7�`���0w��C<l4yp��Gd�y�i��C�D�8���C�f������&��(e(b��!�|��S3V�G��4"�`4��X0,o��`͂��/hĴ_f3BY�Q�Ix����&^���|�@�, ��ɇm8���a�An��c��&�AF����R3�ޠm���p���׆�dj��0�j�	S�0˯`��_����-]C�*��	}����y�����b�FA�9C�G�	|�D�̛��B���a��?�e�?9��[�-��y��62/�Rk#��Ca�U���CMF�
:�M�ғ���,���v���C�m�v8�W{�0������6��s4�)��-8|�\�w�N��������(������v�V(/)AXX���,L^��Z�Kj�w�v�d���.���!"3~!�Ȏ�¤�l,�0;�0����S0�8�!>01�A��02�D@H"�K�(=����o�q���Dnk�e\I�>g#7��f	�0Kjc���FiN��IBaJ%�]!���
�S�%J_N�!J�Ĩ��(���7��*������*q?�@�s �)�������HWi��gs$<�FA/��[����5�_�d�M�؈�udaɃP�����/�di�&��K����&��}�a�kX����T/*ڮ��t�_���ǘ����ո���U��k^sI��Am#�IH���.��Ŵ����'���l��2���e�W�E�/�;�#������U���O��fA�C��p&�I�H��4��j���Bg7��Uߺu[7��-Փĝ���a}�V7���[^��<ŷ��&	Z8��a�I]~��~�!zKd���Y�%�1���5\�t�{G�&���I���]|�{>ڻ�m���3�s�\�p=�o[�es�c�,�^���
1�'��c�1����Y�I�@��B\]�����c��8y���G�|�wwl��m�U�{�����s0vtZ��>���f465���
�ƍ�G���/p��,X��5��ͯ��_Ǝ��//�Ś�;��Γ)��T������=��_�������{�R��/}����Z�t�QD��,��_!\}��]���Bu:��f"�f"�����%r}�`	�W4���)��k�.��:��(�@X^�r����0UkU@�d�J5F�߆y�>%J��#V2	A�U����	j=��_^Ca�0�=���+��0��ض�}���Y���j!v:R<>y\_�4^�&�	bi_*�1p��BU�r|v�!>>�%FL��ykV�
�>|�y��	Ĥ��ըMs�l�}`<1܈�l�8b���S� �3������Rd��������s����O���kx���X��N,��!r�~�)(4�{�j0�'Q_�'"6�A�a��ӓ7��'ؾ� n=z�S�İM������&L���^���� �	�N,����PN8���,\�C��խ�2~�A����'��8|�8>=����O��DvM;!���Z^��B��c&�Nx�<���,����������������#,]�w}�K��a����MDu�h<{�O�Fxf��<����?$�����FdԤ�Y
��7'0=��"�j"*�7U�KjY�B7p��U7k�܏�Ĝ�8,$�Yp��8����7!�Ǳ���+�D�_&1L���4��A~9�0AL�g
�mT[�
8�2���!�oH�i�9���};��3��? �]I�_���ڶ�:�૯�}BU��!z�b�2] �r]M#�5�P7���"wݠG[t�68\n���0���9��%^N������W�K�b�m$�����̘��0f��(�H��X%O�f�e�j�f�kmm�>��p�����4K���ǀ�/��7�x��K���m.�� fL@&rL�b�Z�5�>��cgPUW�U����.��U+0~|'�}Q�����X8�z`�U8p�
�&/�;��)���ڬڤ�]�2a��7[�W�א�4`Ig)f6�cEG1V��cNY<r�<anj�A�������7�u;�L8�T����Ό�MB;�F��$'���� �͓Zq�ʠD�d���&r��ab�� VAV"U%���2?0N��#I��'4�M0��c�t1����?Nռn�d;�uYV�g�[ncJ`�s&���b����f����\�?��J��?����ra�#�퓆�"�|r�W��>�Xz�������F:5"�%2b��o� �L����͝��ѵ�In���>���jb8]�a�D`AK�<tNkn����/,�E��{	P�&H�4��+��!~��3?�/�cM�.Z��# &��T�`U(�E^�F���0b8�o�piU#b�6�Yr]�@_�z7Ä�`X?�{�p�$���]5��Fj���%_����_$_��`X���G��`���c
�_���>�Ϗ�P�p�6+u`�&,�ӊ�S�aZg\��S��pf����\����طu�����	��t���#�/���3mV�X�u��a��w�m�v�{�=;q�/^���;�r�*L�<�G�#?���CQVVI�aǎ��}�1�?���S������dDD�c���t�	6m� E��DPr�x�f|y�>||�f,���O���'X�y'��[ᝐ��,�Xʕѩd��������rD�E氹�'��ʈӒq��Xw��8-���ß��#>=�: }��Մ��%��x&-݄髷`!6��7v�:L^��.��ɻ�#c�t��\O ���	��1��ۆ/n}�Ͼ����8�B0j�l\������M�ޏ?Ƨ�/cȨ)�M.W5!œ���
Á�p0!�?|>�p���˨��>���?Ga}*�����#��j%���P4��+c�pˀ�P�N �g�-}*��"�ᰲy��(�SFLN-&�^�O??��o�{���X�j
�[�Z6\9�7��5��q�°�&��N��Or��>������/���?���W�9uZG�a	/��<�[�c��݈ʮf�A��˶������'���%~6�>�'����O���+��1b�s;}�?;�[����U�'�x��۸�����#m�[�5L<����Q�|������i3I��������v�H����q��EdT���*�x����İJ�cj`I�~-	i'lA�H��K\"	�Ժ�,ԌV��6	L�p�N�[��A���9�8��U<����V�M��=��^��1�k�߃�Y�Vn�s �V�������+���" w�j/,��c�6�B�N5}���j�vXzt�Xu���B!�ǰ�>|���AX�a5�4�3�`sN%��z���1L������{���!�ݺMt H+3�aCK�cm�5�#=G��#7���k�0�4B5��KH�:��e����6R�?���w2�����aQ1�BnA��3��i����8;!�NHH� c3F&!1�#s�Y����.�$�Xȵ���o���a�l��/��^����1�5�;J��� �������%�7����`�[�T��o-�_/���ON�x�Ti�%!iE\Zv��%5�Ms#���,n�.�`��j�����9��f�C1��1���&J�pPL�Us��K�n�ϒ�"��T>�X�"�Ƃ�,�zd}Y�i���/��|�&��=�TWjo�`��O#<���,����U�I��˯`���.v{İ��z��z������0��`��DF��A7êv�;�	���pw������JӪ���x��㠟�wa��wax�����k�o�ҥ+�v�n÷n�­۷�0,~��AW�=��U3���_��O~�aB�'��'�W!��ᛗ��a��p�ۯ`��]K	�%�.��e�1o�PL_����0iT!&�)���,�Y�w7L�٣[�՝��}�S�:�'?܋�'(����4���x���^~��EF~>��0f�̚� KV��ҕk8���uU=3��U�ֶNL���Ϸ��/��pq����8��]|����;�1�Q�0e1�]����s�'(*����������[�)<�{��<��(�m^�J��_���6d��Av�"�TME�B�h]zư/q�_4	�q�KmDA�t�=z����w���>�
=��g�p���p������Z2��!*=2ڙ�No�'����|�5[v�|hʈ�����­G����8y�2v�I%up���ax21=���
Áy�G�3"�n�����w�;�������1f�t$d� 9?S��Þ�����1m�;I�Fp��D��;����� YSV>���b9�Q�9�oi��=�q��<��'�ݴ��p	�DpV��o���yp�°�W:�����dħ�aւ�q��\�� ��=���W�d�2,Z��=Q#�:z��#��B����v�+�&�nqep˅o\!}"Qʋ�g'���Sg0b�Xħ�">%�99<.�������G
֦<�;��pZ�来T��.a��
�Ai�����M{�컿a��P�ЂچVĥe��'I����z=�\��M"��ad;^�\B��\��r8�W��?f�p�!lM�ԞǨvb+�+�~z	��*U,� xe*�+羊a_���Ǳ[B=/.�]�Um�s`��,M#�}� \bIPن�2���1,M$+z�z����mxB��>�c؆���D�n��m�
q��wG�/埁ab���j�G�w��Pσ⟁�W��k��_��R��k�B]�bU;��%V�sRslJ8�a�=�����%^�-����AVݯ�P*�����~�8�-��6�� 2r�)�!#J�#6,89e�ZsG����x�";� #ǌE��1hi�y���n���ETT,�Z���&�~0r�1�3]���o���F�<}a��G3�e`��*��(ļ��X6�Kۊ0�<	�!��0S����v���+�����!�ީjxlS��L�+�*�J�
"�	.����	�h"�Uʙ2>W��hT���N�x1,�I _0�PNym1��$�z��	(a�����.R1�G��	_3��į&>�0���� �x���7��[�N<��_����)P�~n6���T�E�E����%�.��?�}�r�`BXa����+fԀ,<f�p�r�p�wc8�f�D�|�����K�U���İ܈��pE7��N�gX�J���ã0��c�╫�~��^���n�1|��Cw��c�;��������㧯����Ǐ�a�ߗQ��/!�������o��ţx�:�;�>��Lb���سu��3����y-�=���<ьo�Ÿ9�=��Vu�ġ�q���>D����q������o�����������������wo�_�z������?��X:y�+(R�����X;j������p�D��_nn
����=�����l�}�]��Π�}Bb��>a�|t��_��+������ش����(F�X M\�°ux&�B�y�)�]|O��NoGV�<�t�F�9-�bXS0>D�4���JM�xb�.��0�MhJ�n@�X�É%X�� �<�	_�|��?��-۰l�v�߸�?x_���n��N��}!RÜ?���d��W�Hx$�aҢw���x�������k�1S�*?�����k��4����������
��!����P��������������x�����/�DN���GO�U"�ы�q���7����_�hh2�o�gûp��d0��)�м!�+�@@l,A���"�Z��N~��cI�(DgEXn+"��"��20o4��Aİ�_������T$f�c��u���i��r�?��m(�,��/�<��[�����9:FJ�N	)�!�!]CZr�K�TJz�4�IA�"5������s�p�y������GI��f<"��gN�z�rzLsS���~'�	�̥�#���5��E�G�s|O�%�ps;����Z]����f��2ɓj{��^��Rܘ�P8c�������C5w?���F��:̱f�F5}��,Yi8��= R��l�b~�a��'�m�c� X��1O�I*Yz���}���]���;��J�$s& ��a��&ܤ*�A���l�i�ip���58$�6ȇ:����d���n�7s�C�z%ܡ**,��%��������i��*��о�6o@z`؋d�(�A�*�ٺ���j^��~�'(�	ψ�����}}h�ZÇ��MS�yK����QH��|�r�������q��Q$��4�0��K|�VG�f�Ѝ����aJ@���?)�K(Iw��G�H��*��b�*E;�� ��Fz�h�,��;wył�%Öf����� h*������U�|R�4�㠡ڀ_Z�x"�<�A�Fd/v��3?����{a��Jm�V o�1PEË́�B���he+����F��֛_;ںӼ�*�;��{��b4�m;�{ �Ӏ�Q#�>_K��I�����
nm�tXפ��	�/&�oA�So�?s0�x���U��!MP��Xx>����Т.�`z�f��<����1��]��Mu�M3b^�c~x����Jo��{�"�������Y�p���.�����?���;{��%��/�p�������A�8�mF���&SHk��Snz��ٛ�p�H�"��4=���(+.́�X	w'+��A�Ѫ%{)3�2*�6{�!���^)��w/ۅ���A'Zj���h�9Y]��k"�i󥧷с;(�ǻ��c~D;<��	x��F誘��p����D�!c'����-�\�TA�=9;u:k����k��\�@m�vc��c���9�7�]C|ǟ^���iD��4������Z��5��Sɳ�QR��R��}4X��F��-�bw2d���ܟ	S��Iv��4���E�AIoA��Ϳ��?j��W5Rߦg�"���߾rDxsE!�Q��5���n���Z�C!�MNrf�Ԫ�ȃDT���U�2g��WM�����O2x��#7l Q� �R?�>�͜�y�`(�g�b�_����Q@4�^Rd���L3hV���"�W8^���$w�3;3Z!'	
戙�['Ҝ���n5�@��
H�r&��ʇ�y! ��
�Kv��5��ĉ��3��F��@�Є�����)89�>_�$g�uI�$Jm�ͥ����Q)����8R�R���6�� �>�Q@���&��U���2�&���Uk��2O��Q��42c~��_b�� 㿃W�e��p�Y��H��3����3�5D��y���
��s%�����Z#��3�4B�?S�a��H��O7�O6�!S����F$��@���%��Ã��YT��^ߵ��l�N�!�\��R�|=ɹSB�G�a*�w�)�~�(ۿ�x���DV!m?��������9ъX(&�.�е�jZ|1��������!��P6�7"N���|��w!?c#�Q̷G���������M��ڙ}��uNX+��m���C�G1�"W�j��g&��~+�|9�$1����(a$g����S��J"8� .G��wQ���a��	�Ӎ���2?W��E`�X-�N �*�����iN�)'���PJ��h��U�Ǜ��ܝ��K��)� �Fa��"��z�qS�IL����z4���-
^3�p���Օ�>��7��ޛ1ִ����:���_��z�	��o��˾e��\�8A�>x�q�L� �����1c�g41��i����כ�$s<5�M���[��	Q���1C��\x1���EP�ٰ݉7)4�@��L�=qb=2�J�	O|��4��|� ��pc�՝\��C!j
���d4$f[Z��G�UUMȾ�Sn�6�'Z�Y�+�RN��l&����-2;AX��l~���뻮/��W(U�:�إ��m`E)cc��Es��O���lS������^���4�����
�N���o�θF G���N����l�//ٜ���c�J$���p�y�i��h�S�m�H���g�(�P�&�Y�L�^�S�|�;Ԧ]z�n2yC��uk�
Q:�M=�9�kb+��w�\_]9�޲ �/���i�]�7&�ċ]�s&I=So����U�(�}����9���~�� !I�k�3ʑG=�)~��X�/w,�N�] �����~D������9g?�L�����K~r����֕�w�#���dG5J���f(]��,W+�����%d��V�ûUQ�^"����$�w���Y��ȍ>o�J2>�FG��~K������k�&M����6��l�4�-F�r*�qƗ}*�z��g#�")#�y#K\��4�|��yv��P��� ʋ���_Ml�w���Є�ڟ�w�L��jS���'+�Ѯ�XX��/�ɕ�K���s�uT#��Y��Q&/�-j�~�'n`�k���}C*��;փb�����)�W��B%�ES����m�)O�d���&U}�U��N�Jn4(�3��2��O��j�/�����DՍ�u-Ll��5c12%q��� O�~\*?�c�{�`����գ�����-������}P�5��=(��@��~!��0�~�#�8�
]�s���f��<�g̳�a����3V"j�Iڼ|]((���8�r��6/�S^;c�MA�ȸ�v��W�Ι��T�8k'��}��_���g��nJ�D����u�`}��G$�O�9���U*��f�y�y�	0�{����mc��y#�,$��>�t�+���4�M�[��S=s�h���u��V�.���P��\4W+N�P8����䯥 �P6EK����������p_~���8-YN�ˡ�-��JS%�8a�pz�]y�d��Wg-�¼� ;U����-�}� 3�{p��/7��W��c����2+G���^K�<���}�Z�	�Z�54ma_x�'�Z)��R������`��\�W�ɹ�/Z)�G�m�W�]��ʁ��\���M��o���6�����F����}����ژ���v�RE�L����(���sf��5yr�t.�\DZ�Q:ef���cI��E`�e�g��$�N��E������$n||��������i�
5-���Zx�/`7�	5yP���-w�%�n��$�y�Ł�뎆� {v������� @���8Tr��e��"�u���n@@�^��=s'�
�TA!夿3g�U�|��PF�Q��^���~t��d4��:I����z_ƴ�d:����:@W����^"M�#�	-�=�9�H��?���d��/_x�����:��n鋰a��W�ĩ����6܄<R�ޝ�{l�]�;��⟐�����>��P.E)�(U���5?�9�m��O��������'�o ^�X)5�Ǯ �)H?AJ�	���7G��{Ɠdq���!|��K��ӮۏVſ9�S�.��&��=~��bpZ"
�N�<�j[h�٨~c9�`��T��2R��
-8���O���>�� ?�8m�Ӡt��!�_�E�9���,}��1���aOS�`��L�~ǁ���,����)�z�\E�-	쬡�i@��4���K��%/�~PK;ڙlj<�Q�$����l^%������q�/���`��sZ������������'ݢ�J<�rJ���A6|S�Ƕ;�f��VK;�C��}ub�ʃ�D�]��pi���]�W��x$��BiQ��jJ�
8��Dg�|Y�Ƒ���Nɲ��w����^����������������D��GX�L�,��(sm�����PG5~��(���~�np3�7N�M�?@gDI�z7���(S�������)�p`D���e��Z!��s���`.��sqٽiT��W�8(O�8(*�N���1��p�jQa:�Ε���3Fye�.T���%�i����k����ܺ��&�=:��>@]�l Py��h|��@a�qq������D�*gc~Z+\S�����?g�}���Ƽ!$%�"p9�kv�	�793��ĳ߿ 4 76�c�3RAY�a	I�ŰX�Ɏ�*Xw�Z��]�=��/
_Fe.������]�"�)�y�8�b�0�68�Qٵ�3_%|������R��s7�nW��;2-"�ћ���N;�1s�w�;�</zȜ�v;�Z8c��{$�9�GK��6��k)nU?��L���g�$����P�zz�f�u�����'LGSp�^��5G�ȼ�"�31��/O�Јb�tB�k�Vc�JQ��:�F���+�m����#�ɡ���gk"�+JT��4��\��*w�+B\qH`�N����r�}����)�g6���ˣ�ys+�W�wȎ��y�&'���.Z��c9�uŌz _�(љ� ���Ի��}B���9���>�&���35͗]�;XY����a����#�v��H�8J�-��O�l��pv���B��p�!��#���<([��Gh��`�t��ZaŲf�G*E��3�d�I߁f}������Y���]�:pe��V��88�jm5���2��-0��$?�G�s$��~#փ�ȗI��;����`��Ύ�D�9�,�ypk��K�C��}�_(yW�w��6��{KO�i�h���#-,)�]k;s(SD卨���'�� �W<�(Jk;y��Y
Ё�4a̴aݰ�
�}x����g�S��7�F��?ѝ�깜��MkL R7�S��f.��AБ�Cӷ)W��g��+��Vl��	��7<JE�|S	���~x�_~�P���T�%����Gq�g��L(;Q���B�(���Pԉ���)�� ���6s$�3��m��wΌ�>ZSi�ծ�|�S����t��w�c%������EZ��]����+��Jn�&ռ��J��4g�E)gk�	�2I���;r>.E1�����o�����.�U:���Z/Y����[3C��;���E[]?3����}�|�Ò��x������J������1�I�إ	�̺�{ᱱ�&<ۯ�~��bۯ�#y����A?0�=Eu#y��HL�Ȥ�`�%�ʉ���)��ш�.po��aN����\�=��$��|��+�����<n�#Z���Q��s�"�����D��s���Uyo�� �qT�m�N�P靸���kN3Mm��{�~�j�j�c�?-��g�"i�yӛ�gܞj����G��s�+��]ps�N��y�~n�uo�|{s���.Nn�5v��l,2������{#�e�n�U����}o7�I��̑y\���m����\����J.��f�8$�5��yFP<�#���T*R�Vg�
�z{ko;h%H��РW)�}�3Ӄ&�T�j�P�5UC��6�G^`�w��ҡ��s�U�̦,�#�Ȳ�R&RB��-�V�p�:%�}ˮ45=�N�n�d?c���0v<����y�"p�ׁZ�f|;=xD����_����-�����P���L�Q��+W����2L�� r�;�Ռ�p����*����0�E�y���fU�>��~���i%�#p�-����H��n��H�t�!+��I|!#\jvhv�$A�f����͟-X-E�{N��9Wj�?S��s���Z�@Fj�Cd>�Q��p �c_��z�T��9�Lw�u��A��v���C���S�1�������	�uH�;J��P���`��
�I�_G>\Y�}�`�Xq[�`8(��W��ީ��8����m���q�S���&��d�<Iz������_�T��X�'}6I@�dp�=c+� '0��&�xO��	D(���8h<M����hi�P(��it�'-�O�u�e�GK:�}�ɬ��t�-^�fKG9���&GR�V��-M� ��h홶v���1������T��0�����F�JQBo' fxak�XS:*,SW��R�&:���f���*)�
�M9���|�W�TH��X#��Q�]~)\�����D]������N�?�f�~ޑ�&�Il>�����!f9���-U=#��Gbȴ�̵g��8����?%��Z�?��8����bD�ǌ��e}�GAl����$-���8>���[M��*�Wb�ӧ4�@~�8l����c���P���9���>޽�� }���+�7�+��NiB����%�6�F3�z��iRDo�퓻�N,hgL��ƣ�Ts�e����M��z�'v�k�.�.rx�� p9�_���[fs*��TԤ���741�y�BۑI P�28���+���{w6�~��9��z�; :'����SPҨ���,��$.�]���9�DSC�>^�3J��<,Q>���Sg���^�|
�����
��
����b��+��Wi��՟������aڴ�#~\i���[�ibqF!2��N�ny�e��28� ������r�[LG+Kם=ZSg�ϋ�U���L����ǽ�ג�HE�{d3��t̰���{S�e�X�oO�5?7d����ٛ�5Hm�dq^O�w���%��a� ��a�$����.�a\��	��o?i<	�^��ѣ������){�4��D�<��@�l��S
 gc;N�X`�*9�!�h�f�k)��5x�_@@�1G���b��Oץv>)�h��b��H(�
}��u�8~��b�&F����Vq�㲗6��牌ـ��O��8���.��*X��v*�vW��0ϴy�a�\���l�5o?x�[���[�b����Mj�5�k�jm�ɮt}�};3�.��;v�ɢK�JNS��b�_񽤾�S\1�� W��g�T%�m��w�.n��* "LA�(U��p�pP���ȃ�j�O ԯQ��ih曉���ԋ�z�)���X�B��4�P����"���&� �<#�|��=|d�*7�P+S-�T��r"X-��O����)�A2y�B�y�fC$ �1�!4w��HBH�:sA�*!�6}�H���ߖ܆�>Q`uA�ѥ& �[~}%�ϙ�s�R���� RW���2a@��{�f�Fd�?2�֘�k�')sE�r<��u��Ca����g���;=��]�
�M����1o次w{-=������C���	���xB�����O����̻��##9�s�uVs%�hLm�8GM_�G!���%*Z� ᝪ��?��'D��^�1���C#!��oې�:O#)�iAo�$$�&���Z��z%��AѣEG/@��Yx	�d�Sr����y��5y�N�p�f��1��m�P�,?)I��D	ڔL ��W�Պ�&��,kLR�g���e�%���ZC�����a��DDx�c�}�孽����M��&�;��7sө~�/�U@��ӱr�t/�oo��8ޠ��q���ǺԠ���!��9�Y�z��������ZQ�������D���ZE�N^Oǉ��HہE��2���BGe?�N�2^ꍁ���/�����
x���6�I���ۀdI��6��`Pn���tp3���(J�x\��;�����L�����/C����i2���و����R�S ��ȜU.�0	�"Ǳ͟��ƙP��L;�01�9���p�֧
3�,Jr��8�~Ʉv��P��!��1xLyk�4]	�V��3�B{Ts$O�1�m��3M��Y���Vd���E�z�˨��{-s�B(�l�������ʯ���Cc��E,���}t�M�5Y�sd��S}�֒�g�wټ`-��9���J�A����]�Z$�?�b�ihB/�X�m�.���0����Y���Fd����J?16�ܗ���}u�~�{>���A�s)����b�y��ʚ(�G��چ��,�K�D���*��Z��H��x�Yh9I��n��'�w�2�w}���;ڻ��ٌtY��K���w|�R�7k^o^���0����UM�Rz�1]Y�}�u�6�W ��b�&���|���}{�ǅ���;�q*α�C���2}�������?�[�!P)'t�&��E`�Z��^��`eC6o)a��Qa�Um�� �ua�:)p�BV�5��냏]Ő�%4�9�2���n��`�+S��2�e����n�"n�/5q>�^�lw<;=ٟ��8��DX�k��AG�yv�G���C����Ԥm���N]�UU<]/wIp� 4��u�R��<,"F��"2��]��#[����r��}��ylrV����ǎKζ�E:/�$��*$~�I�DH4tx���xt�B#��]R$:ݛ`��t[V)�������͈��d��s���O�pW�=ٿ���+�Om�#٦�|�G��}�l������t)o��ko���暝�$�M���IF�EjV�Q&W�_BŬ�bo<�_�y�<o�c�~�Rԝ����\jI��h�6�;���������n����p?���ֿ�{)���
~g2�<c��L�a٩�	�&.� �F<���	���H�k��s���V�4�i!��2-&G<�Er;�|&�k���*|����	�FR��i<�LV�����p��cLݭUn�E��	K<PT�{���VeV�l@$+^��I*���ޗ�͈�{
3��<%oj��8a�M�#�b�^=��(���mg�eVN
S=�����R᪷5Q� ��iQSa}����;�JG<�_��Lm��fY6�W���y�:����r��X��m�$��'���>#1f��=��h�Y|����&��׽�3<���n�O����O
;��7�Kg�r5�$ {�������e�\r�ǚ+4O�2��z��=���2�]
���6��΁z;�A-��CV�r���s�Wϖ�o���+�PQ,�RN��W��~�� ��])hIQTŋ3�)�r7I�������ٱ���h�)D] ��,���2��$�%Ǥ����?���0�,��q0��U7%�d����P.Q��O�WF=e���N�c������Y'Y��N\YD����v�P��d�+-1��"Ǐ-�秥�J�E��j�L�&��o1�!8&�QP8�*hF����ꩀەkDw\?ֿ��ԉ�.��'�G��� q����F��U�,t��E����o/���bHb�4�q��o���m5��Q��r�Y���4���|p+;{[�3�tj0����� �h��|=R��D������l3�w��RG��Y�f"-�8a�m��|�ڶ�F���,�[�QX�޹��;�%����(-�Br��������6���.&����V,�/ˋ{Qt�4�S6�1U�Yat-�bo�'�哦���Y�N�G���"��7��O��M��D�ci�֐	�+�cx���L��0�Z��U�l?�rp����W�W��u(+$sb�P�|�}w9E@�P�w������́&R9�ʾc�����A���g@i�m��B��^S��^wa�kg�k����ٳkw�S�MӅ�����P�����:�-�I��;����^$~SDe�p���|�0xve��`M�lE�4�R�B@Qӣci���������]?���g�U|�v��ׇA�z@�iO9h���Y����C�q W�n2A�ʲi�8��gg�]įm)!7,u`q�������^`1]o�2�g*�g`�ⅇ�ׄso�}�E7-:px�d��v�:f�M�U��{�hVf����?=ٖ����1.��l&�?
��U��E#zG�k��j���$�5�<n�5�fAL5�T%�K��:���(DAl����ُ��lLd,�F�'Ƈ�D�{1���Tz��}�$��}j�,�/M����;��Kn����,ä޶*�pS#n�˴p/�6w�]_I<��7c�T�=hGs���P��{�b("�S��;�	p%�8�5�C*V�>���٫绯|��J�ܰ�C�����9�W�?�%v#[���7T�'��3�����iT�V�?���B#0G�W8A��c#��x����E�����Ӭ[l��2/r��}����)�w6O'���`i�j�`L�� 晢횾J/��<k ��K�(Xo`ͣ�m���u|��ꊀuru������bS�)�e[��M.Xө��0�A���>���ۓ�H!N�!j�-w>��]���/Sqk���ދJ����]?�B�ej�VNc��]�q���U<F~��K��?H�������/��2�&��M#��o��e­��p}j�~ǽ�c�+�|��hi��4ny��J�W���vD��D|_�-5ؘ�45R���c9]q�6��/��Է���܅�;�;ܴ�S���7	.�i�JĹzq��g�&�+��Td�h����ɻs�lx!4�.�uA��:ҋd�|>�9�,���4��{��̡>'�ܶxlv�w�7�z]�/���M��(����9T�_7F? ��Ȑ@v��uϸ�=~�UI��7�W���GP�X@�<\m�*�#u�Y��vgm±��0y��7���U5��_s�ک�7{��`��3���ߛ���R'�1).�u1h�Qhf�/Ӿ�l�9;:pk���X��3���!��fs���v�����Π��#���V���6R��Ɂ��p�J����9�˧����E21�i���t,RvQ��}x��*g1�1]OH*_�/�r��Z�#Ʈ�K1z��x��'�(�4npQ;���Byо̘��D��٧<�r�p.�c��9/�o#o�Wf��aX[8��f�����4_�Xª�m�)r�Զ���Zy!��{]�E,����Ǒ���?�?Ee�2��ֿ�#�݂>w�I4t�����r�8��;"�0�@�<��n��QϹ�ѱ��z��R7��p��Q�t�ơ>I������I�Hi���k
[T��(B���^F+������NV�⢊n �M�����Bb���t��od�A��N�P����gMI�/��F���3.�?x���?�3�⑂�ܚ,��k�R9G�I�UM��܃�����b@5�ՐoWN�b�� ���:S�R�v�p�?�·��&��;9d>���D|��PW��.F?���@^�lm+*�1�Uq��w v9{�C�������TL �󯈪ϧ�RQo�����BV!w�V����{��X���Ul�I.W"�-{�'�񲑧0vUpzd ���44�|$O�Ÿu��8���[�h���h���{���t�.�O|�r�&2���8�>yCf%�?��BٙE��ҽH"0>K�&-�M��(�<0��Ж�|��!��	P�}�Lֆ\����U%�:���LMd��� ���4��P�U�%9M���9��v�pV	5[�	^����Z6�E����&���?�sg�D�Z��&Jb������$���4aK�w����/���(��q��'�q��1�m�H����=e��D�������w�N��=k�C�g�F��[YjO����\Ȥ��K��V{��j�w��K7��؜Ӣe6��b=1��7{�4Z13n4w�=RS絟�Q��&hqJ'���J�.���_8�+b	K��`�����/�������{���L�3-�/J�������)�b���\?~�/�R�;�N��f�jM=_�%H��YS�%�1��m��ں���`�z�eDQ�RL'H��
�}b�2w�ݘ�c�X�Al]�~y.�^�SV�|�u�]��p��\��X����ڴ�p\͉�<i �z�}3J���(dU����k��6�v��j��O�m�Zy$��ߋ�m���|��s�����Iܑ�5ف� u�_���#���y��D�xa��� �4�l�����׼f��)6W\�_��&6���^���xWd52(4-�3�HC:b�Yiw�++�T)I��&�+�8��D ����]����Ȋ��[���X
;Կ�<�."`*^*J����2C{�J��b��G4�\�M�,�s
w����g	͇�Y���5x׋�o��D��\�QT������k��z/�K��7�	�C�F΋�0����b7�ĥ�7:J�;��0F'.�z�vT�%�MOY sv��⯕E~`�ߑ�6]� �pn�w���� ;.6��1K�1x�o ���?�@��La�h_�1�* �¼R�t��Ř'fJ>��ɧ���őᷤ��>�U�]���ջGm?���P���`yӽ�ݎ���_��˛��O��y���n��$�K�Hx��ʩ�b��P#��ڪN硟�~@J_�O���|Sl�X� H4Cg���,�A��̞Ԓ��V����|��;�V�	D�\���p$vWr�a�#�lnd����6��+�?�8Xp�}�V:�ϫx_nȠ$&*=\,�)ܳ3�
�'bs]���:S�^�j4���p~ ��/�0�o]�h��r>o�X����ӑ'ֲ��+�Vx|E���;^r�W�d8����w2(�b\���^ܻ�e��{:x`ȂB2��=�
!�2E����B�􉼉!��i��+rY����T��[�����r1��Q�� d����(?�Vl@�b%;��f�Y�Ⲷ:��� �O�� �~������Q^�F3��C�e
��������u�tl�K[C�"�yzT��9)E�uh"!g����mA+�su-@r�֎�ŲS=. 0{	�]�x��:�"?���<E)<[�N�Xz��!��P���"9��z*~������&f�m��܂�Qi���ű~��E�)�i6z�知9��~3�gd��,�yuR8�GH�_����t�3ʍ)\���\�'�J!�ӧ�F}E2�j$�f��ڊ0�e�#7�Y3[�㟇��W�s��Q�r5�3K|MNZ�U�>U�[둕L� M����\60�􈬁L�V穟�3W�3���
��$
oM_�W5�T<#%�?Ы�&=��~�y�&�F1����3*�c��Ce҇���yY��1� ���8�t_D����?��˴�X-�)����j�}�3��i�/���ֵ��N��]I�)���Ӷ0���4&v2��~�D�ʼ��9�����G�u�-ٌ�(H/�8M��	;����d�s�-�=V�,R�^��H�:^kP�Z�2�F��g.Ν:��U�ڢ�f,@AmR�3~��
;�!���J��
Z9�~�"�9H��_�).�5�[�j%b+����*�^J: X��^�SM���۪�(��
A:\�\�%c���
��f��^���yy��MoC.9��yǆ��ok<W�4P�)���wl_�߷���	8�@�j���N&��4����{&���q!)N��d{��^b�������W��_"�q�b��
'���PT��x�I��L@���Q�t�su��T���C�jq��sL=��=�k�$�Y�8h�3���5�-���➓�iM�_����5�
��=Z�m�&ᨥ���\6����L&5��3f@p�J��hK6��/5��;�?2������)�pv��q�0ڔ4n?()8Dm,�nR�4���s��}���*%.��[+�o��0{�"x8ޏَ���v�o"+ǒR�?#[Iϛ7jw�E�|�w�֌++�F��:��*�=�s���Z(w�˶C��\���#џ�6���U��T��==}}�ƃ�G��l>�5�X��,�
YY/��X�������֋?�B��o�鲗�1���TJʳ��<�k�   �+��kK�޼��
Yu_���h5��mq,���d���5�e�(u�֮(�z�꾲oͰvj�P T��71(��������B���e����+�Malq��K�{�f��^*��>-�N�s��4�o5Q�ZN�w�au4�Q*�b>�T��e��Ӏ�7W�������r�|ǻH�j���p�q}�z0�n���a<�����py!�U(|U�?����F&|�ÔH�����<f��E�˂`ѷ�EA(���@m����9C/��q��2q�"�"�ru��t��5a<v6���Jz��؀K���x�g6�'��7L�_aW�?���
!{�H�A��o�3bbkt�&�O��xN	�>��v�&�uG�k���Աd7G�2h��'z*[.��}��ya��h�F�ee����Aߗ�d<�R�D�;E�av��f���rۉ���-Yu�)3���Jy�K{�ϘB�����[$�S��}�./� 0K�o�g~�S��]Iq��g�|��I�E����
y"��v��弮ʚ�����wő����G|H\�%E��
��ۅ�f�j�5vysYk3Z��ݣ$���,��5�I#��	)����
�+�ʺX�E(R�D93�����W�������\2��� �����Z�7p�-�2�+7) ~�H|��e�G�3+r�%�^���-�gU�T����ciz�|�`s!V^A�[g�ON�=�$�m��5�[�|��19�7��M��k�b�>��;>�:�mGv�?x��,'b��%���`MO��Ř��ɷg��♧�
�H�'ݑ_y�C����Қ"�K��0�JK�����~������1�d������XQٱD
�6�O��P]�6o�}3
	%��!n����O�P��G���,\K�zk��.��*��(��(�͌T�ӑ/�TH�'��z��ʎ{��D� ���'#��dșE��/�Κ�Q0��B�;]� 4�>�p_��z"(�c������|�Mt̬�XMA�畠r�sI�ǩ�27L�q�
:Yc;N��o'�����-���g�߉:�(�����W�ˈ2I����ɸ2�<�4��4p�N��4�Eg$���!H�<��[���q�'{����$Xc�o>	�7g��K�]�F�����-q`�[6� h��`z�'���(�T����������}���w�<�7��l��O�>չ0=_-��ɍb�׻6c�����uk3�=�$��0����
�N=���9A���z.��/��W'����
7���F�$�&\�����J>B;a\TZ�/��� ��u�ٲh^�55���H�Ǩk�/����G�K!Gh�D�Zz$�d@1�+���w���ռU9�s��z���_�>��ebB������8�.Iw�Qx������pW(Y�;P���/E�I�<��}�M�&$'3^I�*o�|�ӵ&^��2����PL-5�2�EPx�n �Ҷi��1�G�!ւ�(�On�S�q<��u��:E��wk��E���+��j�3l\ �dZJ� 
�� =��)h��_Y�
/������ϊ6�q%G$+��o��ޣ�=�����FrU?���˦⑐z?K�Z�p_θx�����ngg,�\�ڂ�r��'�E���g�o�������R��z�CF��
: ��<4�.�����������8𺪥r�C�������b�?�3�����Ҽ	l���u��W�z#iry���a�݃��&?��_�q�U W�����3����L�k+{[*;
���|U�l���4�A��/%��[J>�e��5�;��Jô�E�t(	�d`_�#��������KwZ�r4����x�؁R�~j�K��g"qFq�nr� ��w���=TVd�Y�&tf��1sD'˘P#�wC!��(-����{g�V��H�O�vo��s;L��p�'TQ�h��ڶ8@��~EO]�$"�᯶l�Ũ3(�/f�Z��O�6�#s�!�NIMz�q[5��")o��I��\�5�u�šW)����v��%� ��ڵ9�ԑ���u�4��T�	o�w$�; ��q��?$ԯ,M�^�b���m\x�▭~���J&���
�	���~��Y�p!_��� X�g��>�J�ަ���?�Hr���t���Ͽ\���R�r�mJa�{l�g	�!� t5|$�4Ѝ���d��\�>�)�H���
�t������`���{�s4�8�6�+���{�t�盒����k6���Jܖ��ߑ���E"3ˁL�*.�j`i�ۨ�+�	�l�S���y��(�6��ua�	�D���8��̋Q�K	�IN��>N^���Dh`
Jt?�nJ�p��+f���+���y��ð��a���rk�*�F�q��i��T:�|�y�f����&�b�Ұ���"��ן8H���)���i�bƭ.�X�4��P�s�[�v��؄9C\2��S���7woy�������'�$B�((��X�GD쿅jF_��*�e�����r�a\� ԟz'ط9\��k����9+=�]�[\��kt���HI)J�Ja�K�t��C�	)i"��� ��������=���/�s�9���Ʒ� Y��K�arg>�x*_�	��!��D�/��ox��/'U��R�N�_��A\X�-J�<8���=�>5�#2g~�Sm`N�`d"$h�a��ca�� YTO�� ��85vnۆ�1߭]���+�g1����<�pG:�8�8:\��8<��	�;�&~6�Y�F�r�)o�1��/[�r����n�	��}7��3���77#�6�+]��5��d�u���&��Կ-&YM��
���椥�}�HgH��wc7`��І��5�!�Jl�h����	� �,�c	���7X
�<t�d[�%�ͯ|04�����^Ό�Ź���	���PZ(���B�)�(�x萿â�1��3�I���t���oh/7��Rp��f�%�q�26xC�=�w3C��	R�u�~ǯ�b��!am��,�7t����A�bydU����I����@�
��տap�E,L�x^5�vb�g�S��Qv��o�KK͟x\��{N������[����,�+�(v�ló�?f�� 3�ږ��Z��|6�O���3WA>ݫ�M��;/��1n�WS����o�:>1l�VP����+�D�Ϫ���Q��X�M��
�+�z����
��B;�1�J\��th� ��?����),���XHȉy�Y��q岧���zn���P������)����7\���S���[>Iӈ!����_�l�F�e:Vy���Ăp�n8��5�m��zo_29��b1x�M�:���{�*a_h���1�b��&ܑk�7G�/ᨪ�RWJ|3�,jɣhc~_K8�
D]�kd�y�$Е؜¬~��w�N�ٝ{�R��"^�D��?��`�B,'�-�ྻ���l=�@���N��н���|������tF�R�]��)��N�I�g?��s|h�3��եr����va�&���\��/�<��Z�/_���H����%k��,��+Y�����V�4!'
r�����Kl�egJ���^���Dn�۞������Q, Heb5��E��'ߨ�S1�����P"���Xm�
.�*�!
�㯥��/��t��+�aޚZ��Q��g�Td5VO��v	j�.��\�4��.������4�V��MPؐ
2*�(K�������`T�q��x�00�5p��u�������/T!~y��ځI��?�_�:V��}v�➼|�E6�u�|�������R�⫝f�|ʧ��T+���ɸÑ�$O���� Ħq\���V�2X�:�|�P�/_�w��d-fW��<�#�~��?�����&�&�p�������Y�k�V_�E��\���:X�v��\�Q���A�j��$�����+;$;��֝=C5�+�T5J�=p"H��5�~'��B\��X���S~�	<�z�o��4�E?���5�tr��&S�:��>���Z� �����t]��KأL4���P3��xEa`�����֮�_�k�=�3pO����xb���������~���9�~4�֩�{E-�-?�9�Q�èO���q+uaר���H�}������I�(��`�"49V��?A���\��)��Ī\�%2#a�����'~�����n���$&���mp�/r�K?��+�!��Ŷ������[�y΀��wY�����#��DS�Vc����H="��"�����r��Ӷ��"}�w�Eg�iz�Ͳ�S���z�s����R��M���sU�m�\]��C�.#{���=
��U,��E��z�g�-$������2�t�Noﵯ��2\�,�2�'lw��d���c}fK�g(Q�������~�vMbekIS�+2���P��԰���I��/��nl�Ľ�GS3@��*'���j] �s���4���R�k�R��I�5����/��˿hX4QT3CE[��Ox�Ȇ=���\m"�_���+��Q�v��M�o���"��RO�}Do{i-@m���<X�D� ���7�i�R��5�w��k�r�2-�
��<;�	)�w��P�j�m|�<�LLt?���9vO��-<r�P���W�#�3*-�D�a.����?�] &�Y�g"���N�L�-�[&�1*��qh���w/�М"����
�� Ɠݩ����4�o����"����H��~�_8^%0�n������Aל�WG���~1ͧ��	.߫M6n�3ʍ!����i�������\\$`�}{��mW90Lgr~��1ğ���.n뾠��}�T`���'F�E�d<�q^�~1@��Y׭uc����ͿyR��|Ca"%/��a��h�ο���Q	�ƶZ����Q�سA~Ϛ^\���o��-^9�Q�Ɵz�xH��=�_��~(��gv��r��.�gv�>���kkH�i�A'}9}��-���>8�����Pw�-����x<-O������%cp��]{��FA�-�5�p���
����.�- ¯�=�{i{�畄f��3�޶+�Q���'�Q�֑��կF�&�?��kk
D��p�ʉ�i3�ڪ��q���e�t>�$0n�pm@3}������v
�i,j��¶�Իm��x���_��+l��H��;��$��EȠ��Ha^uƇ��@;�ʤ�߸���P�'}�`��(�.k>��1��<r���޿��:���6�F�R;�F	�t��]�P��**�"W�ͥ��3>��k���*�H�-E]lw��j���B֌I�b�6���'�n^i��>��R�`̈́���!b�??��M�n��4H��.��ǰO��v1E"�3�����)�,&��rj D,>y�2웾O�"/H���7��RD��'0�6�]^���u���/�w����e��0��E�6�B-�b�S5�E�6I�SS�+�tM�g�W~�S��aڙ��U���	�ߚz�>��;��x�t��p?q��3iw���?�7�r0�/'	;<�P���dٞ�a��
�<���8ݝG+_z/u�Mn8�rV�������v�	#%£]^\6��')1�p��c��7~S�53MV)w���"�F��K�%-#������{�Ѐ@�+&on���[޼�!�nlv���%�:�X<f2���K�ᗼ�(H�c��š8��MXT�4y����ґ�^*�jt0��}��ox�Xx#����cT6�U���T�d���k��������ɚ�Crt�|�$�f�h���L*)�"�1s�m?�wa .O�f�uV�@F2�K�zϖ��@:�Ro5�[/�č�)[�K{��`&���A����	����*F\�G���ѝ�q�,|��B(,PH�^y��ZG�v�(�[" ���;�Z�"ڲŗ|�7>=]U��e���B��ݜT˾aj/����r�@뇄6O&���8�=ƈų��jc{�w��"����c�V�d�����h+C36'�/3s�
xd�`O�I.�x�,��H���xe �c����s�WKO�M��S�z����@�%�p/�_����}�e�;���W��������CUO5ڋ�qg����2�x\�ε���`�#�_�L��/�ܵ/�vpW��;���$�Q����Zm'�Re��N{�><�t3�e����_�D|�w�_=�3A��g�$�4�	���s�J_1`����g�"�-���長a�2Pj�g�收^5*gC�� ��5@�V�i���!T���\\	�?lt-�F�N�iPP��|�aP	�b��Xޟd�ɉ!��|��*����甠��+vQ�ο���X*5�+�]��H_b�X��Xl��\i�|w2p�X��%��<�5����i�毾� d���\�#�%j�>���Zo`^Wy���R�/��7������Vz�ߥ��.o�Ə�x�I�
ǉ��@G[Cy�=t8b�K��_�������9���Aw1�H�l���Z�uk<("ƃ�?&
����v�_���Y�.�i���hG��;@/��`��8?j� 4@�S�!u��B����0}]���l[��	@��0�y(O&��_S����.O�{������TUѲV��v�@�Q�2�1�]y?P���#�GSu��#p/ݼ!�d^x�� ?v+�J���eu���n��g������-��W䁔QB�wq�5d���X�E������)1�X�#����f?/gR�m�2��g�U:)��/��,5�r�)>�,|�̡�{q�2�s���4�l��/��of��G^�Bngi3oɆۮɆC.w�/��,[X��8�+�{� �'��C0��ơ}S�)f>�2���tT��__�����,�wC$$�J�,|��)➇껰s�%C:$8�BG>ݦ���L"\��btI�F��]��'e�k�����Y�]����U�{Wߏ�eq^��g� ;��+��7�X�b�.V����F�J�/�W�B��~ok���3 �a#��f��if��S���cCTї��w.ڙ�B����5���ŏ�oڊ��}i��	��:�l�����%-��L�n���o���W�hѯ7�� ���Q�.���������!�_���Z�����#}^�7s%��]�R������T�5F�^��F¿�[����7j�i�[@Z���9���Q�_���y���:�t��A�~i#<f�A<S�U�U�+�� �B���y��:U$=Qe��6\�l��Y��j��"�.Ξ���[��!@V��3��dzl��Y��C�"��//���(Bҳ?Ԏ]"<9�s`7s��$K2�Vv[{��~�W��4<�(���@�����g`_a`���ﾖ5�H���CH�v�<���H��� Wh�'���S�)�4VR;��`�#J�n����+�������!��6�x'�mU�p���)5���Gb��Yp���7E�-bauZ8�.��Qc�)�C�)>%�k���$�T1 [�Bl[0����A�ҫ'��׼9Eh�����T��=����t޺D��ݗu�Ra�5x}�cHq�o��eD����2[���>ŏ�*U�W �Q��q��-���G(��5I����	�O�����.���ү�K6����u���(�ް��6�:T�_��bM��ݫd'z=�H����#t���#t���)J�N_�sQ�JJY|ttFF��i�r覞��b~�:�yd��(���f/9�3�-d�>���|lD�)PO^��=N�=�bC����^�@�4��X5\R���H/����oB��S�w���l�����@��^��;Pp�n�?�w�����?U)+�T�qc���va?�~U؜�^Y����ܪC���,�w����#�?j�p���3��;E6[i�9y�pH�"��9�L���+�A���\+��Hs�J���CB$����0���<U�r>�+%������@��뙷SoHZt��I-?ؐ�hD��/��;7��Ѩ��k�&�&db�hr����'�� ]
1 ��a=��0�ew3�M)�5���D�z�97���JN��&�|���2�I��P	�xo��j庲Z$�~F��S�z�jטc�0Z�%]��<�@��/L�܊R�Q�c�!� ���vK�*!�VA�������a��ӕ̏	�kg%g+OL��g7����-Ȁu5�� ��A�ݿ��·n0袮���+ ՋK��h!�[n�-�?�ō����lYM���I?*�����[�5��6�!������Y�M*����~"e+�����Q�n��wX��T���f. _��� ���O��%���hM�~Z��/��9�4d��}Dye�!>o�Ʀ��_����/��V=T�~{+�C'إ���ˣG���@�T)�8���΅,E��u�<�Se{����<�A�O����"C��SHS�]���'^���D΄�¹�u,{;��<���RR֋����)6%���'���ʇ�7������D�*��>��Rj�Ʀ�Q˚$�����VN��E!*��qB��j�:I�Ć9��G���@�����$M��C�4E�/ ��/e��>�s0�ǚ��j%���o�w���7�ē�ݘ?��^��pG�\�`fT����iY��L������A��"���ܰnF�Ǥ�2�Jch�11�岉A�^�p�9J�eb��2Єlr�cs}�ǝ�$�Ï?�$)��!D�i���&�2�A��V��f5�pϒ5�2� �J7����(�\����m�Ix��:3���5
�O!Y���|F��`����	��z���/�5���f�����k��/c��$aa�o/3s�Re2K���,$)�#�^�|��R�p�(���Y�x�$Eg��x�^�g�ŷ�� -�N<�X�k������W@lX|�T �2����ab6��T���JD_І!�
����BL���T������@���qk��9���W�G?'q������������w�(�~�c*��s~��;�%��ʥ��%.�y��SE�Ey�v|T���e�$����*.钍b&uw�����J2C���2Zq|z�Ž%�O
��Q��&��]/a����;����8�E妵`�����M����>e>(ϸwG������c_]ר�n$�)|JS�П���CŪ'*?�:����6��IQY��������}���P���s�6��7>���cߐ���#�Q:Ɣ�MI�d�*���0�J�΍>_B�����&���dY�{��C�+%�+8~��\�
!���`z��/a}ߡ{e�C��ϭ�/Z�GG�@#����>%�A�0\���~;���}='�,/_�f]�j?���;Vn���N�!3���#�?Lph�Ό���<g�==�P��=Z��/�װ�0P%֙��wL��u�adX�ڎ��!���C��U��,-H:.�p�fk��0�P�ft�
���˱K�aF�����^�9tǭ��Ӧ�v�Ԁ����i�֐�(�����K�2;߽72�=5Z������Џ񍯍�wq[���%���tч�vyJR4��7*���f��R�~�v	ȊR��q����9 ��>]�'�w4NΥ��2 \�o��{]�\��-��6�/kM��=��Cz�LmJ���g$��Z�&(̶?-6�^l��ޯ���9�=�d��q�ܢ;�30���E�Υj>װ.��f�{���礣���
��G��pT��(���א(t@h�=H"�4AtN���n�+2G���$�=�R��}n{�����J��T���?��+�"���2�zѓܲ��F]��3�ڏ���ՠ��f��_Hp��@'�ć�|��#�~u����yv��G�t.@���:�}x����Z+��d?իq�������������aP�g���w���U[k
��@g���N�rs/��6�yQ�������}7�,3�Ax�&o/O%�����>���B�&��=n-������tQb�|]���F���<�O�8ʄ�[�ɾ����*��r5�|���4���9Y���ĈqYi�y}�Rd�^��#��V��">U$��u�]��?g���nFG!h��(G���^��t�m�j�ԙ1U
١w�*9����Ȟ���#�;����
�6�\�L��<�e��B�B ��`�V�W�-.����gVW���M'0_cQ��md5�Ȫ
�9��'���������j�i�8�~dR������������G-0�B�2Vש��r�*�@�q�]��Vw$�sB��7�!w�-��¹�����1��Y��r�hg�]��/���a`MS��~8��W���R��i|Wڋ��8��+�����Ѭ���\Z:E��Uw��{Y�eF��}�����|e���n[���"�5����R�9���`�k��T�@Yta
ky:�� OLK2��\�n���qQ��?�����;*G�"��A^����z�b�Ne��:��j�|�Q�Ґ���2�uF�:�
��0jRc����f',un�0O'�ʺ[f�(�rS�CУ�G$3��{���l�w��fe4�5QH��f���(F�z����������<�Z��wYv !�[��J�4:�Ҍ%��&��cHǎ[���Y��>)�� (%8	�#�K{�T:�I��|׿ۦ��,�HV��,�>��f��C!F�VSvI�*�{�Q�}��4
�QV4^�M��'���G0.̃i���ә4�Y�:v	]-�+��y�O߿J�O@�Q<DO%+~���0U�a�\E!�4"x���a��S˺Q�Y�
^�,�cKE`��v;ٖ��{�x�h�kc/#`��b�+>�E�u�q:J'J�	��ׯ_Q�>��';ӑY��+'��m���mlS�j@B����+�JKO�i���H���M�'��z�읎�t���hnd��ϑ��m�m�����K]�Nveof;޳u�c�wl��pPe��;��b�M�<�O�t��)��U]��E�f	�in��gr��/dέ����/I�)��L�:9j��՟3F���H�?`_A�H�Й����/+6Y/�W�/����"��Nô��갲�>�9 ���X���D6����ᢧ�_���G��3����Xr���?��k����x!JQ��%R��G����Д�#�����2@5R�/��#���tU�x�Xf�T��z5�糊��w�@5��c�����߶(O���vp��Z��Qu��Wt�]w���;�Y�c��������̞�<nH�IW�/4M�HN�Z1M�D-��\�����n3b��*��r���ś��a�6SSӸ���<<7$<��R�7�Wb�11|�º�qr��\Q�m����_rgEτ/��	��rΖ}M)u�n�����T-2m`� [b+���FD>�C�I(������_��v0��)���M���ܷ��>��X�Z�0ƻ|��X�F�p��W3iz��������E@>�o�?)�_���F�.����,�����G����I��6�Y5��[��1tX��N�>�v������1x�lb-=�� ܇��Ȅ!6(�F9�b�"&�W�'~P#�$���ߦ��	F3V��>�(�@�'x��_e��F�3�p�.��c�܌� O"�Ԝ��|�vّy�b?.����^I�$��*3����;gQ2 :�Gm�E6�M#h=�!��CP�U���J��8F;��x2kp�w�j��J���"�M8C\$ep�|���D� ��~��8\Pz�M�]��w��7����Hh���'v����Ǔ���G)��ب%�5(�'��N�*�='a�2��D�N7+h�E X|�w���g��͖b�������������.�Y���V����@�!��h����Ix��Gu�_A]�iĿe�U{����J��ǈP�<lKGR^T<D�a����Bs��Y�%(O5��OT��u�R�<_1[�	����ۗt=ٞ�0�/���"-�I���A�@���N��r�׿�W�|�P�~�φ���H�+�@g�~�� �b��:�h���S���q��$��x�O6$�e�dt�� ��殷�LaP�>����È10���g�N�G-ŘR�п�P˧��|�!. ҷw�N>�,$�E���Uu#�w��� ���QϚTŌ>�0g_	�V*Ȉ�IX!XZ��j��1��W;g%���)��~D�^�jMX��`�F��C1�>U�����ֆK?�{s�s䍊�.ĀD`�hDe4@;�(�4��W@�s���(��c�9F���҉�)�Ԗ)��tρ:��G��,�~ES�	���q�&�6�3����^IF�RH�^��2 	(�ҞR?��k1�'B�8��ϨP��C�a�7�jv��T����S0"_u�CZ����&_%����Ϛ���t�)�$�ϑ�ٛd�Hp��^D�?g���2��C���븢B�}�*�<�1��ə�F[+�͉��\�\Eensz.	�
�N�"�ئqg�f~xTtt��'�/-��'����.�&��co�.��)��oϥ��{�_�c�7$�
q�Il�X,�����t#���4�������E��4f��v�d*���7/X;#f�m]#�;\A�|3�q����YA��`�G~�C7�g��X��&����2t�J>��^j��Q�D�0m��}��$��K&����C|�k��Fc@��Ӎ����`Utc�[3ۛ�?ʋ�O�o�6�3C ��ɛ�������(pQi;�s��K��imH�/�G$V8�^LIK/���7�$�C̩~Q���(O��R�;沣��hВ0o�B���v&V����_�+��+(^2!{qũ��=-c��@>�Z-_ �;;uE]�����
���4�u��P�8N5�Ѿ[@W�]����UKo`T�aS���æ�r��i�v ��o�SV�����y&�?M�L��>f~�\�]ƒ��u��7`�r�v\uL��S������뗐|9 ۟��Gk>{�{3���A��e��	T�s=�h"?I�{7���Ɲ�?��3����T&v����� @�7�����Oc��Q�QB��oأn)��*&y�,�����Ж��#�@������t��7[_F$wj�im�J<�J��k
{1RY�������o.�З�� CN�Y$ݡ���nҁG#v��m{{�Ȋ�o�)�N��F4�|���G�e��YB��"���L�-���G4����/�A��x�[�T�w�Q��A+aI���4{�Lkq�_�y�+����;�j*Vq#��T�a��iVxl!H5��h��+����8����X�J�Hu���:�n(+�v��Bd��*��R S��@o$�Љ���^'�{?�?�~�����l���[#�9-��pY��z�;
�b3���.�bz`��_o�"�/�0��K�3�1 ��	�w��H@�g�>�:�>�M{�W���X7����FrB�[?K�|U�b���b���������|�nL�7 �'3�J�ʑz/e�g���IY�^oĲ)���[�ѳ���C� 6���%��{Q�A_2HV��2:t���5)��&3���8�$�����Qs����f����r�?kǖ4�E�tB�1��'�%)�_���V.
����-ks����S��~����ZB�/dh_��*�X��d�:*(������:�����o���'`�=���mj�T�w��A��6�Fkд;�P�:"��;�jV;a�nt��oP�����>��Sk`�;a%�:�"�	?��~�䟩r�`,iAd �xp���'d�9���V��1:�C�_d���Ͱ���<!�(�� Lmmdr�t��j���ğ�
�E5($�6�a?�������޶��K�y�����[U�sR1tv5�ԃei!\āK���xqD���E�~;� Ġ?Pp^X�$�5՝b�� �ډ�%V�~�0����̠��΀[s)$0�҉�c��QOq�bG�9�P�����,�2�j0��q\��M4���8�?%-�?A��]P�u���hd�I�����c��Q����:��Ƽ�])u��B���sza�=�k�C�ŏ�֮�������^��5�ɮjG.c�s�&�w���?��y�ƽp��("�e��x�O�C��.�y)�v'���Mi��T5 mѐ=���Q��n�'����%_vХ@��r�~"�����!Hч����ګ��s�3qݧ��-|�?	�?������N|�:/�%U�SZ)�y�%.�T�i�yV̧y�x	�R?�1Y��>iu��joܺ��՗m��\�䴲E���\�̹M�$���������t/�����p�_�y�\*��К��i�oo���@,�'183����AA�Ϫ�b���U���b����߾�46O9��|ԇA��h�-v�킒���ɺ��V�\ )��!n+s���r���.U��]���Q:�->q�
�~{si� ��ڍ�³w/D�3H��w���H�N�q�f�Ran�#�0�9{�7��Z|�vچ���;�?���t�^lm�,ⶻ#/��w~����F<��=Q{H�}�`*��vup�^�����Z�kQ���B_[+!��1�Lw@��3��I���g]�$�=XF�ǃ7���TiU=��kܷ�ց����[A}Ӈ���뛪��QjNU�D�+j�!K\���W��S�b�]���9�t֜1w&��B����7IW�ީZA����8H������r�-Zv������2q|����ք�)��M�ժ���fLۭ��tZ��u�n��cq⨻{����Z��H����Sg,X�4�ɍ��cR�9�9%TGc�e��G87�~e�ȗ���)���^ǌ,*��D�RH� ����:e�Q���Z%~%��Ȇ�rLsʧ|Y)H5sf�2,8ƃ>r~�'/��c�K��������x�gm�v���VivM���Ի���6O$|�����
o�|�t���B����&T�_�?f5[ ܖ���b�hD�R\�u�å,��~�����z6/Q$Q,�O.B�$2�5�\��x�r�Bu!v�4�aI�q�c��gPA ���X���ś����0_{ƫ����%�����LwY��3�����$�(1$AQn���e��v<�Uj�@�*!��I���-\���ܔg<��R���R�)�qsD5���,H҄A>6�0�����zRҲ���_�Ԏ��>�`�Ｙ�L�ي88`H-������\�PӅK��ɣU��J����[>ؾ2�.r�?xI�[���+�>�5s�?���VH˓!�&�:��L�w�����M&j�t/�/.����Iߎ�#�n��SG�����R\9���{��Ȩ+�JU�^}�㏼���M�*oj�-~\��{�U��h���:Z��{��p�nBӕC�E*r��
r�Q���eCcs�"��̃}i75����%L�Ow�֜��p����H����G�Y��7�}ւ���mސؗ X����}BL
����I�fǾgY�l��j�]eb�/�!3X!���xAѝ,�R�v	dah�ؕ��5��l�wc�>����pR�\����$?\�lR�'�b�<�j�~��Љ�&����6��S�F�\����ϱ�R�e�����ǉ}b�q�km]n<D�[��5pl���3nã9�E��V�#�D���G�"�wu�l�B�'aI4� �Y�f�C�u��:6��{����)�����2q���A������=�K��y�.l|��z`+ok@�E��,�q���l�d3!ű��sտ�Ǒ�b�Yqİ�@Ul������Y[HG��b/�D��<�1�����؍z����Lh�L����>0߽:?h�ɣ�Q�7	�,���ȭ����%��K�/�YW~���N^���]�I�����Ű:2��C�Z��F��F�U�����b��i{���G�&Ke·/�1-ށ�W�Tn �I�>�V�Y��Wq��ai�Y�M��vڝS9�q��eԏ0�O�Z����y�Uo���#8����T�I�Y�[�(W�ĕk�w��� ˲��%��������O �!�k��0+��^��u[���N#���N�#1,=;2���I��H��� ��)��¾����P��V:Wg��ot��(v��Zbz����?�|߆ٔ|ؓX���4�\�Fjm��+���/���r\�d�+���U��g[�~�sJT��K,�C��;��Q"��G��?_��Rq=�y���$S�n����%��/b��pכ� JMQ
W��f2��`���	��s+g���i �6�qÜ]P�:F]�(t��{ƒH��A�/u�7S�x��/��`�Ӊx7+���1��!��I�-��i���H��oC���*uֹ�Yܿ]���Y�u~>�77�߲ȍ�KR����$���>F�Xx�H"�Z�sn�'U���
g�^�����4�e�;�6��A�k�Քd�ܟ+W��%W���o����25�.*^��5�4'8!���i��p�|�P��+~h����J�&�cZ����%~�d�yr�([ŚFwP���%��b����g��n=us�
`�������:��S*>ߵ�p�EG�	���oQ���Yz��x�|�5);#B@i�c�=�&�\ȡ²!e���V��w�Sm���f���'O/"����o�s���2)�+K�%$��n$8��9Ղ�d�Ą��߃�nfT��\.��Խ���I8t����2S��.�&UX3_�m,J����;��﬙<����l�)17??:i��S�\\Z���)��Z���h�õCl�Ν�@�f��e��K�'�&���G&`9&�����f�0��-�P�0�cآ�vԐ�I:؇/�m[�r�,_�⑻j�J_y{h�~N���$��ʊ��e���!)_ޒ9⡓��| ����H��8��V���]�S��$�k#ƥ����R$�r�k�4���ѵ�Ƕ�(��z.�s��.d��	_�0� �4����և	\��7�Vg3�smA��Z)��=���]��P���x��[�����\���*!< �~���@��k�X��CP�9�NQv�[���z�%4#�!���ު�	)H���
:��|�G��w�9�rq���Bhro��	9����8�/+����iekK�C\Q�E��y�j��Ҿ��Y� �#=�����'���:Tų���$o�~"����^���]�ץ<R�[:M=A��k�q)�xz����_ՔH�8�_�:L�i.����J&`h�컿�A�#l�m �f��G�;���K'jJ}͝M�{�?�^1���sWި��� 8��DSWo�ܒ�.�b�����-T��rw���� �)ь��V�0�.�#�C�ӗ�[/�d���p��x�'PA:�H/�O��	���8&�X������%�$�O2A#Rp2%�?�E�|	J��)C���3zFV�n�1�0Q� ��H��S&A�Du_��a�GR1FP&�s��O���>�������
�B�|����_^W���N���2n�ɼL���i&1�G�o���æ[�i�����'�GǊ�T��:q��������f#q��Y��p���%0c���+: �����C������)���k>d�ŜN��G&|-�������S۾>�s�=��2��n���J/����Tl��2?#�`����9 /o��/��������Sn��Ey���a�-����,�;���:����y��E�x�T�5��^��n����G���~�>ů5���������*�f'���_�3�z���/A�?�2�f�I_�o	;B���ջ◘�&���q�x����M�&�~M�[�]��zNW��'=�y��IUx��qU�s�U�۴�7��G|t��,.�� ��P����os7`�+je\��8���sS@qQ�OFv 
����ltKBi��_���L�:~���%�6'�z5~�/�K��Cj�@V
�ܲ���j��@���K���w  0y�y��.V�\u��W�#�?G��u�͟w��{���3����+�]�(����P=+��g��8!��\?���&�8b�<���ŵ�Bua�G�U ��H\xm�����[��ʵ.v`�?�� ��~)�-��9��uYk˺�3p�0���@\�f�4����[���x�Fpo��2�R�ҁ�.���=�x��*�pY��t;5��)�d��u�"�g��,@"0�!�ݎh.���q}���B\�w����s�xb,�������_:��Sd���f�5�ꔿU�p��X�,�N @��e'�ߌ�A׃\�D*͛+��Rh���-���lՠ��6��7U� O�N)Q�
�v��m�M@!����04�?;Z�v�v&�%h���.-EAu��uU9���gֲ�������I����C����[��i����|~��q���ֲI��аr�확�[�s Ք�"}�lk�ʬ����%��3C"ę6�$�6)İ>D�9�w��Ș�kJH@[r��K�nx>���S�>9�t!A�����+-�)�����ɲ�]�B�����N�����G���	���Vz�	ԧJ�W2�D1�-���_E�|�#8�����$8^��p�Y(+��L^�M����#��Y�^`E�vo;=ګ����$���t���7Qw>���A�Քl^̝7e��bN����j&�N�R��� 
���e�v���x�T��K����7�2����<�d̝J�J����=N��O/�N����Y���	��_�Tԧ����z�R >�ԉq<q�yV��R������B'7�,콻�U�6��"���-�	�t�^�z�'��]@���	C�;�?���=xܮ�C�X��*1�+�NE�p`A,�lXiر��}.�X�X��������-*�ip>�桳:�f��w:L=�a�s�h�߰w��{ ��b0n�T̜3OE���E��^X�z-�
J��䎸�D,[���-���3\�пO.�����J��Y����ߌm;v�cg3���9j6oَ��|t�Й��%K���pQQ1��MP.˗�@qA):���IX��"�:v֎p&x��;kV���t�h���$l޼#G��3��A5v&6m�a�Y����Aѹ�����\q�X�q�	�����7{=�����^%B��|A0]c�`���%��Y�'�⾒Ө�d�9��:�j��a�� [��c\
KG?�ZM|���n�4@5�Fp?�l�`�`��n��@/+�f�?cl�U1����M�ۮ�!U��~ջk��DS>�T[K��V�d$�s��x� >���I(D)K��2�SS�vm�mֳ���~����w��Ė-�q��<~�GO�GVql�c� Ð����2�����wp��+��JF9�'/�å[�q��|��6l߂��J4��?Ǚk��q�a�բ�_�3�ϒ���� +ޏ�ph|-y�j�&�ܾ5��%��5x�Sַ�@'�@��	�,Ot��y�G�����>/�+j�Wۧ� ����5��
�	����
 k��2�u��w f��&�<u u�a����*�/a�a��0��wĝ���0��E�ma�Mz����?���eN��a�e���K�b�jlٮY��\��`X,�7����/�� ���C��#|��1�N Vb~�>�^�a�C������`����ھ�O�ţo�*������,,�7C��(W��r	�jZ\&&���2��-sp��Z\��	.�݁�N���Q]��.6����N�&�hi��v�`����hg��m�
A'�(Xz%�%4�QE��.�w�&��l�&W#8�+�3k�Q	��rdW!��N)(���D���
��*�fV�'�J���ٵ����ܞ��냀��/@����&DW'`�A~�(0)u��`D�#�N#ORa�|5��N� L���~1s�ׁ�ȧtB+�/�a_��N�
G����s�2���++��J���!�f�G�Z�|	�A��ʱp��F.�C��/�KbO5�rR�Y�+���ᄋ�c�$��0ٍ ل���P3r1r�)k��3�E�t��[������O���2�`���$��ՁNE� ��?�X��S�U�3��W�It�`8���`�Ԟ�N�ރ���Q�����v/��,�M����MY֔x��5!�:BK֭"J4�<�Y�D��g%�ʊ=4n!��K�oX���N�����s���Ss���c�51!��a��ش~+�,X��x��ѣ�'Μ<�����7�GaQ9��;�5�����v�M0}�l:t�)i���'�`��Ř=k:w�gW���+��Ba+�N������U``�!x���s�.�ݫ�[������"0 �ۈѣ&����-1q�<��{���������1.SY,~�9��Y9:�9���J�:���7��V�o[ð�m� �L��26��؊�;%2�A�(�L��|���y* &�����O`�zx)��4 n�\|?|���kȻ�t����9��G���uR0K)˷�b�O����@����)�$�"�$�X��r�>k��<Ow6,�2K����U�q��g]{��78���?a4����l�r��x��LVq�-="Y����3v��.U�`��\��^�`7V�	�{�t�{��0��=�������G1{�|�ط����u�>��q�I�{U�{Z����-�aX�2�J���\�w������@,�ĸ�!Ri�\=GJ�m~��X�LU�`J@�2��d�����*ݒ���zn##V�*"�v&�Co�`BlЫ��w��;b�t�k�l=ow�1:5��@�f6`����:g��a��6���mZ�p�|��Ka�������,��y���0w�,[���l�W��&_c*0|�0|�W��K.x�/���>!��p�~ ����*�� 6��a�m�������?}W.~�`��=x��f���L�n�l�W�qCK0et��늅3���U�����~i/�\;����c��&�'��o�7����un���	ö�ho.���M��_�A��/�{L��&��Y=��)���}Y���}R��=\���QՄ��A����ʁ)����5/���o��}y»�F!�zB�G#�j�RXױ�'\��������\71��^:��O�%WH��H�[�9�K �x�_�a�r� �*��_ú?���W>IY�ehg	��Ŗ�i(�p��K ���|���p&��#8�&1��k[��[R/���DJ��Ax�r�`�S{j���a�5#�L�M�AHA?eY��s ��'�c\J7^Gr-LXЉd �P,0��g%0,0)��܊�W��R_O��(�a�M��?���0�:�X��re	t&�'��3�AM��GA����3��U6^i�U�?�l[�Жpjb��aX�1�b�����Җ��՞�'"1�]�K���Gd>�#s������F� 15+V���7"08�����;>څ��8;�!40[7mǪ�k���OHm���=p�ˋ�ѽ~�۷����v�-am먢�|��~T�W�C����ŢE�T��.]��S��h$�غ��`mf�Ѐ0�X���́�w�r�<p>�`���;�����m�g��	0�l�N��0t�|~�<B�S�v�p���S@
�	$!9p ;�r�g�-�D�7�l\��`XY����|��&�#�|/�a$1���̤Q$$��9��y��iq��<�R��q':�2�
,+Hn�#,����D[x5�\��x( ˴�4�Ĳ�T���u���;,�r�\(�8*�*�����-��2�s]�\���1TÃr�㴸 �?&Ù�f���@tz"�]��/���S�0n�X��9�c���ۯ����g-�_T*,=���\�w#��FK�pef�A�	���cԴIX�}3���lی2XS}-��Y�+�����;͹���h�'��G(�@^��[�\��j0#��eJ2��@y�� �48D6Q���cF�
k�2s��F�� X��͛aX�$��p����
��
6V�Y�5�p'��9س�u/d�aq��`���x�;��2�b�&��Vi�C�.n :$�O�a��A�;o�υ�N���g#:�uG;yS��Ng=�[�B°X���X�����ҕ�����L������2|��mܽ{�g���p7��x������E�����*��K���o�X�	�?<��i"������m�ӧ���Cj심�S
�5�^%[9Bӏ��o���a�G��r�x~�.���_���{_���ؾ~.��������0j`�."�*���	��3�����e���q��\>���31~d7�gG�����N��7�ۣ#A��-���O��:L}e�4��g"<��y��(��i�o!7�"�DvK���ʡ������a������	�U;�]G"�nb��a��n��e\Q7�ݰ�	�6!]�4��d������Y�$G�c����!�hJ���m�5
�Y���0,j��@(ե`���#ŉ嶵&���b�}��e��澾�a?�a+��,�aӐ
��K#�F��'����^�2��}��.������`�����B*����g6���	�v�Y`�rsٱ��.� >[;VbbY��j@@N���d7"�����!��ຬ�����c+�*�V�QR<��Y�*5��D�H�SV��8����l��WY�|�C�M ��F��I0O�2K$	Ձ.�0�,0܃�PK@������3���W�_f|2d�����X�3?	�D�vf>��d�ag��ȉ�+I�H�CD!C������%�+(~!�H�*����������
;���_�AA!���ADX>\�=�{ô�9l,lU綅�������o��`�����������3&L��y����������8L�>���������Ÿ��Q#|�d�ڪ:lX��5��ᝎ���1����8�}�Ψ��K��$g���k���(��*�^���x��-���y��p�P0lF�aeh�JX`�>�����H�0E�t��`����!X�nn�b��/2�� [h�@d�����A���+�6�����+x�l$yg�Of#����;�|ٸ���?����-���2��5��j]��eJ�J��3?�����&�q(�d��m�y��QS�fI���(��HE3ɕh&̋���'
��,S�Ô��:��6�Y�ϗ�k�R���*bi�8���5<a	I��p�fe�ÿ��|�-�6���i�)X�j�{��<C��������n�+�����&���Æ���Y۠T��lg����p��m?10�wF��&:�%>9|=�F�! ���1��0���
��"�!�DxT
#�*�!��-�$XJ�c�!�XRY �4�+���K�/��H�zd�m,BĔ���$��\o�r�Xf�"�*z)S%B0Yd��Rn�ve�f*a�^�:��B�^$Vj�v~3�:���u�]^ï 1��
�e^�0���`�1� HN"�3	úe��0��
�?��nh5�C�q�7��X�u� ֥o��}��uZ����a�W�_�� �[�EX`��ׯ�a=��_�a=ư�/_@\%�_
�xJ=������������������	�����B�x|�?��j�����\�����P5��>������P���[jɟ��nS�p��1����<���u��l�'��g`Ѭ��4��c
�i�k0gb=N��c��1ذfvn��|��ۈO�,���Xi�����;����-:�x���?[�!0󎇉WL|���k�2�'���1��?�sz�ao#Yx���a�G(��A�K�p��E�5�PUG�6�]�j��CXWB/a7���m"ax©0*��&!�+Sn\3��+qr�0�1���j:�b,$.o�8^-� �!L��aJ�a]���0,�+"�*�yj)!XD��'�4k�A,ԙ6��G�ˇ�����X��D.��e���@�� ���MT-�28Erc��#�+<���@)�:�y�ë˵�Lh�=�8 o0�-BRO�D�p�֌�7+=� ��M�赏(�+A$�����UV�l�'תJA:�I'2��f(����X�+,K"��tu��\��#��G��t����Tj�7��@��'�c�a���V*)'���l)�U~��xt	�&!�:�� vK&(�!��2פn��#`�Y{��U@X�:���q� �6���JG1�-$ Cra�
��b��&�#$��N�Ų�>��5��O������`�(.-�����b�طw?����[>d�|v��y����!�a8~�ּ�>��?�ڱq:h�@>r�G�prr26oތeK��Ԥ�-�0k�,�� *J+�6�;+=�?ڍ%�����fV�2q
>޽9����?�9Y�ػg?�L�s8:�aժq��%�'d��?����?}���'6�Csa�{`�;V�v��hB��ɲ�Q�0�]+�Q�1���A:+��U�B�X/���yv���X6~�s��<��Al���������������|z�	�Y�LbVB�H�O��'@�"6�D�����2�7��rڏ����ڞI��^�$Hz½y<�}嘔:&%�K�/�Km'�s_�_��+�y����*Y�Iy�2z$Ӛܹ��k$�������I3�^�)��������`���z�?�ʍ�u�<��_�g�����ŏ�g'Ρq�d�� ���㚡l(���d�s��|5�������#�f�_�S��v0�X�ع��; v|����'G���)D����;	��հ��!�,��"��D(�q�!������JJn%�-W*�tik>m	�b	�28�� �i}ކ�1��A6��K����s{Mo�!p�,�\n!Ӕ�uXd.��ZE�J!�k������#�d"+G"��j��G]�?�Ȇ�� � ��dP�\���L��+���7 ��Kk4�Þ�K� X���E��V냷���,�p&:�W�5��R���a�!�c�aHf�A7t 5�϶j�\�^¢��"9�17�p��$�΄��I��%�:�ף�H��0��0�|�*lش/]V�.}M��-���I������p[�e�jЍd��s�k��@���H`�A3O�������P� ?���?�x��|��E/��_d�+�֠o��}�Al�������'�'�On��[x������,{��N-0���^����c���؉{׎�Ⱦu�h��غv���NQ���t��؁Ř4�3��b�����XK ^O ޵�]ܻj����Ы�^��x�Nh��
��\�������kڻD��[,~o�0	k�~x3$q�O�EHV"��!� G��)��rB0�H
������Q#��d�j��Ԫ��	�� Rkpq���"C���N%8OQ
��m%r���`EV�i.,�@h0!����7���hs��p�Lsy���Xkş���E���-2�g��7��H���`�b>
��������\��Pf�B݋0,@,��, ]b	��B���^��M�K���̾�"�z4�1U#�}�?�ĕ(�P��ZeU��b!�T�
�X�:kq��U�� ;+P�e�F��
K�8Kُ�+1���+�+�X��°X��S���XZ�?4�f��%6���h�abO��nı�.� ]b
�@��#�m��a�ůU`X,���5��N:�8��]"�	��pHW�;�'�% ~��=p���
�7oC\b
b�╏��N#95������_}u˗����b�bq��)\����~���hj�B��\����o��O�݈˗�BFF�����sg�bŲe���@TD��݇c��!;#f�j��3'�`���pvp&k�ml۲Q�Ѱ��ô�3q���6t:u2CFz.N�8��{?Chh,�����-]�|`��86�`���+�0�ǆ�D(�Ct��WA�50�{�
S�
�)�]@m��;+~�9K��;q�	ȉe�.��ŊH>��W���c���%�#�oT���EU�Z�JZ*j�I�������*��T���|Tg&��%�R����H�-T��ŲRL*ZK[^�jڌ�ά���>m��ʗ�d��.lH4�N��:&���Џ�)�0䗋β�?��ɁY`!,M���a��=���;���I:����]񋗏p���8r�0�m܂^M#���86�h�*�Upn3[�i0Mp"$�fc��8}��,��@t��CHL��a���PL��w}�̊F����e%�3�aqyP�� Gj����Y	�H���H�i��l��u���D�pP��+Ɉ���4�`4߲Mż�iul����cH�u��'�?�I�Mz_���;�9���{,��\g��L@8�e�ި�dCJ�Qy��oye�#��1�r�.|�os��
�_��0�\3�߰O�`�*��T�p+��Q�'�i��x�����1�Z~��7�k��y��^aQ��$_�3l�< �
�{(�IcF��)C�������Ûՠ�҉N�a-�į��^� �������[���f���O�۟�b~��{��]��{W���|w���
�޺h��y���}��� N�:�on~IIzN��o�e^���cB�@2!��g�B�z�}������.���6/��3{�}6���-�O��1�0~X�������1~H�����	�X2g ֮�`�}ⵓ��i����{5+{[G��_��[o��������`���x�.�8��>��O�gL�d5<��w�֙����
�'��)]	����Z�*���Ո �`$"�&PA����0�_D�T��g ��l�l�"��|�u����y\�.n���}f"�j�*	Ǖc�!�K�.'�Vh0,��e-0����@k�M��%0�/�`Xs�hk~#�|*&Û�a^�;�e�l�fd���:����
xŉ�p��a��Z��	.%�U�;���NBހH�1>yx�c� ��wrWزps$�����?2Ӏ��pJ��iP���������k
 K�4bq��e�$��e���*�hv�=չH��ҡ�)���
�ĤC̛`X@Js�0X�yn.˰3�NF[�A\�����w�18.aYpN��w<0e�2�8s	�,GC�h4�?�D}
	���:`�X����j�8{[���_d�+���U!W__��'�'���������ff��1c���Æ�s��HKű#G�� O7O,��H�������U8��Q,Y�A��ņ6��3H'(��_���u=q��}�\��6�pv������l+�0��'��?	�)��JF�%@����sK:ǿ��u�Z��jh̨�Tפ�JN	�
��3��fj>�%�����[I�"��H��T>W��60�;n�3aY$�,��a�R~����b��>w�ؔ~L9�7aE�r
zvij��I�o��o�v�ńp����k6\�~,]2�,��b��~��,˙�������7�zO¡��c���p��BqY�]8���^��QC���(�����;�^����#8�^�-sa����5AF�4a9���	��]�w̼���>a�%ǒ0��AP^�'�BE��0�J P�����w��3J�&��������(7�`Q�+�^�EH!�k��K��nIP�h���a^�k�q� �c�9%�D�-��˴>/��~fJ��"SJ�4�����/W`؂�/��y���>
r���R�wϞ�5i��|[�{'�*P,��@���Nð��t�3����y�U�V0�Ax'���pK���~�Kk�u�0t!��K����	Æm%������l'y�e�Kr�R��SBtd9e��r,�uav)
z�âe+�ߨ��t� �!.w��"6aMm��0,a־'�|� ��'���Ӈw�۸�2�_9����ܩC8yt/��G�����O����q`��ط�jvo}����';Wc���-�2�r�ڪi��رi>ڴ�7,e�q����|xSs�P�a]m��z�a�"��<�����c�B\= ��8�=[���5�0nHF,���ݰ`Z#f��za��~X>w0�[2���R0����X�x8�Oj��aU(+L�������᝷;㝎�x��o�����?޲�B;;_���v>1pI��G��3�08�'��;�n�0�Q�����|+킲aĖ!�����3�'��G#�bӱ�&�F��QǨ�Ɉ.�FM'�Ma:��WI�c*g �j:�ϑ�����$Ml�������O�aJ�a�{D��S_b	�&@,��K���aq�a��*�0�NKg���i*��X�!� N,�=X1GFT�Չ͜��=!�>�������|�
6(��#�7�	���&x%u�-[���TOB��]!���F�V*�dha�j0�r�P�l !T:��EU�h��82j\D��p��M@W���_�.�!�ld��P�H,}O6�"	��,�e�wN�?a=�W�s
�)fZ����we��SB.�aϕ�=WR6L�a�tx������W8&�Z��{>Eo�gYU5�M��}�~��3g���VV�6}���e�pw�P#��rsf������X�D`` ����?���#���ame	ss3L�2	��y9������DlݼӧL���?�C�`�|��#�6V������=�`�x6�0)������D'1�����QSU�S'�a���03���W :u����YX�`�
�XyF�1 ��IpπsD�c��� Xb;;�kԡN,�|G��F�u3SK�����H�0,�{W6��ĊKXt����j>���*V`��{��D�#��\�՘�T��L�f���X�_R0�i��과�NR��(1c"��|���O߆i#)�2�EWk0���m�.�U*�1:���ϩ��|�ce^���3?�/�l��x��w��|�㣏��1s�\��"�9�>}���o��ᘽ�=��4�6 ���ꋁ%�F�ܳ�<��l0��0���/����;�q�+���ox6�}��_�BPL&�����W���e�U�E�/ao�j����<��.���<9�\'� u���(�TgMi�dx�%�=�]dZ����k�l���g�?y��������׷�J2m$���T�R�]B1���B=?u�Q�������cY�rL��|�pOkP�;��@��z@ ��u�p;�l��`c�uw	����eJ_�%
7�K�Yx�@�ɏ�a8�0����������`X���2l��Ӝ��d����o��H�O|�m�Ӎ`�e�Ûp��W
�%������Q�M��K1a��3�x��zL=����ٓo���Mܽy�����.��{Wq���_���Ӈp��g*=��>�:�1N|�>߿	���@���]�c������,�۵[�ϡf+m�`6���kE����X�|�,����'`��p��<�E�K�� ��W�X�ŕB�f�@��g7	�ߵ��Gw������a�4�[6�{b`C.�,���0or?�p#�F̟�������声b�0L��C��!���p��IǷѹSg��l�w�ؠ��:�z���L}Б��O$�݃a����l����'$�J�Op
�)��L�G�  � �%L�DpZ7x%0��Ip���a�)�Ċш+�鑈*����#p&ULEx�h��S�f �z����iH���T�z
���U�GPL������-
�����f ����a�u	O3���X���>��T��S�1���+&��K�����i��{\5�ݦ"�|a�VawV^>:/�B|��qM�-�Oy�	���W<`.
��)�D��^1	�c��;���	��Ch�X���k'�oˊCB�9S��O>�	��Vkq�%��D���@�X�%�T,b��5����(~%��q�3zB�κ���%�t� ����u
�x���\+�0�Ʌ�S|���Í��J�s#عŖ�5Zb7�-*n�yp
ˆgt�ӫ����	p�Ő�S1g�rĦ������yX�b9z��+�Z���@,X�Q�0�b���D,\�ݺ�������>|�r�PQ#BB��~�<x ��akm�^={`�E��HS��s�_�Fx�{"�?M��0i�d$�&�����9m�w����'ܜ�0�i0&s�x°���	���/A�npv�BdT"�������:��7�=!���Hع�3(����W�9Q�@o%b��'m��y��/Z"8S."�����-��/�[��U���ni�K,���15
�����yB�� pA7��+�U�H�X\4��V86X}5X�$�%:���@���LtpUpJ��ѭ�zx7�˕��u�z���ռ�O���Xw���u��$c�+��f]��z}Z˟�N��l�������#<|�.\��o��������W.��W��gx�g`�����9����ĕ�Q^�|n�J`�����KL ��*�ڏN���;��=��d�n��i�>�/.���k�`����(��[������A9���yg^�)e���˂�Y�Cq[��I�	�[��t|��9kQ)�)>�R�%���u�e��PR�&�T�|_#Y��5H���C���eb�[�u_b�!��8�ݐ|�R���W��5�5�\9-�ݞ0* ,�X��=柝 +kq�X���E� �/~S�.z���0܏0��ľx˿�0�M�"�q��9�ax �R���G�����G�"~z_'}[�����-���AXD6%���a���a%���s��g��wx�>�C �A]�����/�0��� .~�)Ξ܋��vQ;q��=8|`�m������k��Rj��'�c�E�x�h1>�h9��X����峰s�*\�x/�0 �V2����0|S����+�b����M��գ8�g5֯����G��g���`d�2�ۓ L �9������t�p,_8+����9�1bp1�xTG"=�.�����F�o㝎��N�hgj����0�wG'+'���
�^������?£�����d*E)<&�Y��K+FXBcsW���2x""��#��pd�Cb� �	1}�����ܾ�/����ȭ�����/�G�B�G%�,K�фޱ
���NDD�xJ�I���4�����0�I�5c~�u�����.�u�&�0��m�&��VM�O�tNOG �8�r�x=�Y�)�;�	�
�	�����ራ$� +�wJ���#�iu�LI�������b�z��5���Z�Į�K�G�mf�DQ�ju�R�R ��b�F*X���_�<����&��U`��K�_�d%�\%�g8�^m'�
�ǖPnr.2h��r�<[`X$`U��,�D����󠌰�f�n�a7V��a��l��"��F�z5����VvG]�~�����b�0`� Tw�Ahx<}��������HHJV#ȅGD�W�>((�1���N�-..Q.QQ�\�� 4����l�����9Y�e��ё
�GTd8�ס��^�^�7
�ѻg��������:��* �NvՕՄ�D�":*R�~������M���Sq��mܸ�-��<���?F^Q%��.��pa��3����+�E�ݔ$,���{&�����s�b%��CY�=r�sɨ.|���G$�b;B��C,��a>��:>�n�B���܉��2I��T�;P�|�v"nk[��f�gi�wA,i�I܏��,�D������z;J Î�i>�U<�iP��$f�kbw�G�%�d��ĽC���k2���im^���x�r9^[�rm���e��~�������i�D�#P[�4��>�ϳb���\��kW����o���k7�����o�L_�Au���Aו�	�(��d�v7�?����H�bYF�g���(��������;�=��'|���t3�lBli-̂��P)�s:���a���ώ���X,�)�S�N���x�� [�K_ּ�n�<w����a�e-�s�m%�5��}u��^����N��b�r^޽�/�yIe���Χ��Kr�ֈ�rI�|57y����~\+_�	�](�u:�;���[��p���`8�� ���F"����1�*(�`�Vm���E�}�d=���1��e8���%��K#~J~B~L~��>=����ݡn��7���A���<����ȧ�p��-b��-�Am�,|v`%�w5�z{>��];fc��YJm�O^���b���س�}���4a�&�=����]'������Z�����_�2�t��X�s'v��s�5^9gF��<���ư�%��^X5��?,��ų�b�aX0{ ��3�4`p�<t��!G %�vVo᏿�_x���wo������C�Nx�����VG�ݾ"����S7x����/!��	��@@NAd\Bc�����l��K\�L$ԡk������F$�#6������q�{�FfU?$�#��r�D^�A͒�ܮMJ�݆ ��4�t	��&��j& ���[6���f��aa��A�+��%2�����7`X�]3X�%���ϯ��VO�_�4��L�o�4��?��/0,�M`<�a7���5�tsf��Ax����j' �
a�A\$���DJ�X'n��BX`؏pQ�_��܍ם�[�0)8�	�=&"�|��ƪX��jÜ�	�i� �m(f�(0,��d^�0A�0�A(��lK-�D�Ns��2:��CJ���:9n���K�bUV�
�a��K���>%B��~h��5pg>��UT�cK��J�#��bװL�I��~0v:������- v�tĦf�?,ށ��@j&����?�pJ,�i�HIˀ� ��"����lBrBB""	ұ��� �&$�!6.
����c�����"91�1���Fb������"""�<~XX823���t������S������H���!:2�i��hu�_N  ��IDAT:i���̂��,,��I��a��%X�d6oݎ�_�G��������|4B��Fn@NO��BP^�#}��OŪe��NH^?��Q)w �Q�%�$�CK�2&۝�DV���Sz*I4_���ǰ��`-�$
CM�K"MH�J�(K�����WI�5yf��|oE�9E�疫�7G��'� |$R���D>��k�D�ТA�Q!ZԼ�y��|$,��m^������Hz���D���r�܌%q��7�����A�/�U����(C]�Xl\��Vo����1|�P�=�'����1q�d�Y�[�F�1�a����z�9�,;�/�X���?�Q�46��J�������3|�OY��ӖbĴ�4i.��F"�@bF�����ޅ��,���<W7�#c�]����ܲz��H��KV/8g���.��d�.�̞J����]��E��1��v�댧_�k�SǠ�Y�i"����@1�A��2�����YN���Z��r,`�@�H��Xh����)�P�˶��yL��R�"�,�����2��+�xgÄ��F�z6�7��W UW�md����ߒ�g���1t�aS�p��� _�2��p�!����W)�p�&����ҁ��/�@���Y�E�x��	�?�03~�@�}w��E��o�^ŵKg����őOp��'�^M�&q����!�،/������b��ⓝ+�g�R�ܺ�7�ö�s	���m�Bl|>\5k����;�����*ڄ���|$baIox��b���p��M����n]9��;V��яp��qd��[13��%砺(Յqh����q�X�l
�_2	�����e1���4aδA1�+��(@����L	��}G���..V�CTB�cY9�$���I�i��O�Сñt�
45F�����^����}�P�� �!#Ǣ�� ĥ *9U�1j�B���,߰�������{�D�a��G�q�a�����5��(�ԅ���ӓ�y�4��;��~����Ə�`��/�p���h��N>����GL��t$|�)��Ú�"��6 �@��4��Ô�!�0�¯�a�ր���ﰈy����OX�s�W0<�0<�0L ���\'�+$
��U��>���&��+��o<AX�$�z��!�.�]�J#�~
rz�Dl�h��Pe�R>�`� ��ԝ�S2��<q�Ǘ��SL5�c�* vf^����J'��$�6΄vX`VA'��5Y�&aê��Vce(n,0�ŷXbs��b=�mt�����M
te.=�L��ry�2-�����@��]S��F ]|��%QY��%�P�b�r_��g
�r��V�+�L��KΆWt6�c�X���%4�����j��a��	g�`��G#8*������GpxB	�b���ChD8"cb�1�C]ph�7��� 8))IY�	�bNNN@Rr<"����$ '�l��m�-"2<���d78�<^l\,�;�侾�/\#*:�TlL��Y <J�GD#>.����D���A�������62"��	EjZ2��0y�\��3xyq��D�$����etCHND��t�Rx^oD�5"��D���;�I�%���<��J�/aēp a��	�Z�"_ �pb��"��ϲNM���X,�ZD	Mv�|�YK��A��|�bAsN��Jb	vT�3H����|�tK��V,��C:�5W,��o��c�ƣ��Z`�Vdd�լݭ%ˌ��uҷ}�������_��T��)nD�_�#�T!�l �R*��[�08�E��?�~�� H@���{D:�J{�'�]|�a���S%d��J%���\�����n�0�MC'�$Xe�* �I��O�UP
L���7���&�E��2��Ϝ��ے��uX�d���z36��b+`J�i�|��r�D��3�%]&u1�D����l���7�s4S�95]�Nܷ3%i�H���d��1��m��s�	�3��Ρ�0Q2t�#���;ω���[���X"�H��!�?����P�}�R,���7G�K����\�q�b]�%�fG6D]s���k!����	*7�p��x�:6M�v�C�>iW4�"�g3�t8���T�l%��1�y��+�k,��u��:�!��]�{���U��b�{X���=�n�R�ݐ�~Yh�W`���_�������f�|)�'�(���x��>�ݹ�K����S�r�4�?�C�>¡Ov����[�g+�ډC{%��zՉn��e�rlY��ׯ����x�:l�`9֯^D�]ܬMk����es�n�<|��ܸtR���^<�-Ä�'�	��Sb�������p���صeΞ���9�c�b���=�;a89ɬ��rS���h�Y��V���K�!}1i�P���B��"�U� -)��N���#�`��w�clھ�vmî�wbڴ��ׯ7&M�m[7c˦�`��Y����9�sg�ĕK_��կq������GZvr���n���z_�������p��},{#f.\��g������<��G 1����ջq�ۧ8x�,�}}߽����-����W�ǭ�x��H��b'v#�EPɨf$P�U�}U�`�`5���+0� ���þ�a�.K�4�d�:5��@o%���x�^a��S�W%�ƪ�t���������ܔ
F��'T�R�N�gh���N� <}���V7�'�	=T�K��rx�"*��d��~���k�2z�x��U�  ��E"�`2zLEV�i��"LH���PK��1��jþ���� #�Il�l��z���+&$�'vU�,�M�)jR���Y�!�|��0��u��H��qŽB�X,䲝X������"�� ��" �`��@� ���{�Gf)�8�לAN�oB|�zG'(��$Ï��Qp�D��B����@�h}���T��������2J�����	�������z�e� �d:A�[:��q|).������Ǐy� (8��	��/��y�3����~~�ח��5x���ήN������9\�\�a�0q<N�:���ô�	�m��	k���G��G4B���FS�p6"b��W��Nl�I,먮J�|���K)>��P�)pZu^S>�|��	���V�w�ӑ4j��4?��R�_,�f�`c�`J�CX�_0�I��Jj</�0ե:0�y��;F�Rh)�j�ەT��w�8c)�a�_�_W��q�}��X���j[���b�6�'�X� ���H(S��n��ET`��7�<Ӹ.!��6�)�ssCt	צ�#+$
�|��E�t
�F��l�^����w����¸��Ex��(]�n��6��ׅ2���)	�#�с�T�o^��̳�������#�����.����Do�:Do u���X�x�}���Z��dZ��o#u�� ��|�:r^c��J�v>��P��@���^���?��� �o��B��6�L�N��a�-��U�5Y�<���=�iM�L�`�]p�h��.��0�D�mG�G�}�0tHI�4�p�l:c�5 ~���V��fc������	�v��p����[c���8w�"nܺ�`XE��yK�!@�K`X�� s���0���c����op��\��r7o\Ɨg������K_��s�r�$���.}y�����eܼ|
O��{�����u�4�\=����0=���y1_����q���ڍ/>߃3G?�����I�"�?=¿���p+����ګ0��b)��a��7�p��'*b�y��/�ޏ�`��=e���c1�o%�v/@��Ի��墦8EY1�M�FeA�sҐ���PĄ 2��!^���Cff<fϙ�/N�gG��g�`߁��}�f�~o9�,���+���ի�i�ؾu#V�Z�5���m�p��gl|�e�y�~v ��MCBj�N�����É�W0v�1;�ƽG��-�г�P�K�q�1�����ې_V��Ɓ���i�=t��NƲ5���ş��W7�g�h��� '���� ��~���(��ґ)��$�	��:�&�Ӳm�@�� ���0��,����D>���V<���Q7�5kx$��p_6L}6�`�n+!��7�V�p3�Bp��X�)�ٗ����:X��̿P�@Htǘj�,�����>�b�'�z�e�=�I�
��{�@n�j�7=0��tF uI�@X�TbK��V W�����<7S���N`X,��,ۉ�X�Y�a�G�k�_�W��a��c�KH7�aq���N�y��"�wI��侾�r���U�$Bp|�-�q��D�'��;*��p%�:����v�>p��y��^�P�_
����~��|@ ��K��%��Q�$�r;M�'�j0@���K8n�{����P����G8��5��w8@��|�xa�@o^�<}���&0ls+3t1��.�PSS�+�#?��dnGg�F�a��.�0q	�C@��R����DX{�QL��aC�&x	�:�q�P�
[�{�Y���O�:86���~ùO�fմ���[�$�Mô���V$����Q��v�{܅ e,}�/]��>�]��
*R,$L�k��z6t2�R�:�,���Z �5 �H�7K:�^��MRy�{\�s�3f9#�52�LxnZ'F9��s����&���bn�I�(
�0d�9ф(aҌ`kIEv#9�}�ٸ7�$R���Bxq�.�b��	AV{6�@lP���.����ԑ��`�L�R��K��N�����&�k�&}��s3R'Q8��9v��sx����w�"�������r��4�p	��U	xK������k�~�c�7
q��i�1��|)��nT�Ĳ���LkP,#�i���(S��R��<���I=��դ�p��B�ù��\58�߆a�σa�h��vc`�φa��&tI����
��
8疱��E+Z�$.^��[w�����J÷n��50��0��0��~��ܼu�����%_ĕ��p��<��@*#�=�Ͼ��e������w��]ųo	���d��OϿ��{�p��s�{�<���wj��F�2<3�|zO����_��/i��b�I�������O�x	į�p���������c��%�]�|� vm]�u+ga�q��M8r`#�l]��˦a����6�F�# נ_})j�2Q�����P�G!�iX�"B|��@��8������Ŋ�c�G�p�0|��!&��ٽ;wl��;�w�N�ۻ�Z���GcԈ��5c.�����b����ѫ��]�m�^\�� s	�1I�HH�Ÿ)�q����a;��k�o�(��p/~�_��ac&�W�!����شc/*��ĔY��0|��udV�;8Vm�� ����Ĳ���Ȋ��� ��J��p*���ÚZ|�[ð�t ~����0�e�O`ؿ�	ùy���7�?�+ϷJ�|8��G���	6�Ù��vO����Z��@��8�UX:ѹ�k@t78DT�.��@��ב�������ʍ��8a�Fߴ^���5!�M�e�#ǐpfJĄO�]�S�ܨ
�0aT:��f�FJ�X��e��	�¯��n�'Y�0���0�Ţ-�c�j#��0,!��B.1��E_�~�OV!ٽ�SO .c#��E��/C|Q��+�AEed!��E�jQZ��Y��`*�����8=D���A�ð���	�˴��P�O(V"�i�?�G�}UA	*����*7�ѱ}y,_B�o�'a��~pqw����,��}�v�й����۷c��(,(��o0ܽ�����1p�T�5ŵ��Q�Y�Ȯ胴�ȯ���aHoPQl�$�DC�'��$�])�|>��M:�HLh�@>�K:�z���zq���V)���h��e�F}"�!X�O[Q�|������(k�ؒ�,�o�B벋���5����cۉ��z�xmцk�ѯ���A�rh����A���4R[�	cw	]��7Kbr�S�[���,InPd����ˇt�s����/W.M��BT�����U_�8m�e2d�Et)�crQ�(�5�����#�yK#Y��y/�y�lx�t���%�[�9=f<�9˟fqʒ�H������G��X�q��t�䳓�8^�kd#�g��U,ϓ����y��k1��,5�W|/u�郎���Z��%�le$kJ��I�Q�1q�Q�@�]B����G:�	[��(�����LG�ϱ�6��e��A0�Y�Z\/d�YY-+�����a���o�2�0Z���s��7O5m�^�=`��A���j��1��g�pg°	a�=��v�|v�a��r8�!��/�]��V�R�0�`���#�ƍ�p��[�_���q��F<�B����?������x��6.]�_}u�K�D�xB��Ӌ�����Ve�8q�!���v������%����z����_��+����c���]�~�@	?=��3���R?=RP�����+�k
�z.#��+.b�5X���H?(_a�o�8�W/ƞm�߿qZ�L,�7K��ʅ��v�t����;�C�TbP�J�]�~ue��(@e>�83y���H�RP���P$%�#9)]kJ0z�L�2k׭��}�q`��ٵ۷m®��㓏w+8���~��1�̞��b�䱘I ��qz76`��1<|$��:�S箠����N�@rF���Q߻��;�iy
�Or�����ظ�c��h%�\����j{a΂���%�����j�ɽ"н�8��?w��P�8]�D��BD�x�(	�bV ��aM����'��b®���e�/,@l8/�t»a�z<|*�p�Q�c$��7�����e�A�JJj���I,�'���YQz&� d%��=���ك��W�\%�ڛ�k:2��A�Tf�L�k���0���@q壐�}
���Z>����r,�!+�*����#�0L0�O�aC* .V_�J���"9�����қ]`XF�r'���$�+��c0s�.��p�nރyk7bƲ��4Vl܈�~�Ac���eK�ɑ�8p�(V�[���Z��D�/4ބ\wq- �&��K��#4��q�.B�(���}�L�U"��}�W
�T,Ⱦ�Wo«7��G Z���ׇp�KiVb��Dx�}|�|T�	o/Ox{S����ec؟���z���YY��̻����I�8{����?���o�e�v��و��Tt�������ِ���>؊5�w��#gq���8r�>?s��G�ыY0@�O����O���{���_bC�%J7V����u�SC.�~Ǚ��t,2�3O7�����ۻfq#�S"�L��O�2t��1��R9My˰�J2mPjO%�qv�>nI,X�q~�$_+�ע��)�Kڹ/�#-�;�w�{E��a_c���{%y�}k-_���L�6��J-�ۅd�'�r't�/41��N��i=X&4��>pZ��'nk���mRl���^�́�D�ɵp��ٙ�\gn���JG2�'7Q�&�6r�9I�
��rka��� ��)�&r��{���3���K'EY���7�3S ���rg>n�ݒc��9�\Ա�\�̩�my�x/=�N�{��sr��y�N�Ǒ�Q��>M�u2��<�$�g�|�$"	�K���P��ٲ�yg��,؈3�:��w�i�f���Q��2��4F%���[���?Oͷ� ��]��z�dj0lM�Jꇎ!�a�\t*b#�����j�V]m�1V%YfP�m��y]^"�����,��%� 6
�IC&�����Rd�������0�e��q���o޸�[Q�0�K}��a��	���	���_<�Ͼ�J���w�~�/�Ù3Gp��g���Z���o�o?<!��W�[����_|w�?�a�	����~xDX~��	���R�������~��-5/p��/�O��s�ۆ���'w�b�}�u�5���?X���Q����燸��!�ܼ�`~O����[W��i�0eL?�l�Ř��1jP-���ƀ����ǀ��أ
�TzT�GU���������$��㢃�����|�ބ���)��`���ظ�}j�����»�tӝظafL���c�c�����tfc��?y���3.�����Z�i9Ũ�3=�AC��Je]1u�Bnw{?=�Ϲ�+����S�t�.�_�Mm#����cgQY���(��s7��|�ƭ�^2q�S����- �K}�5�Z�B�B�L�L��I��0����I4	�G�F�WRÕmb4��~%���T,�yA�J,]	M&nY���GA:��(t�&�`����/�Y2+�xЄa�͟�g��X�i�X��ӏ��i��EP.��.Bs�`\�>;��tI p�]�v�'a�+]z��K��ŏО �k`X@\�3$t��<{��U\`X:�	$��Z`؅0�H�`e�wÇ�-�&v8�������N`���xo�&,X�{?;����b��	X��Z|}�&h7�n@Ͼ}/?B)��ېj�
��ہ��?� �l �X�����H@��*�� ��}�â@o��E��1�|�W�6-0���7S//�{z�T:�y�CX��ɴl��	Oww%/w�/0L����c�y�����f&pwwEVV���Y(?��;:p}z5"$(���X�~#���w���X��V�;p�O���ż�;P7p:�r{�&�|>PR��H*x	E����C�ˊ?���XًT��(i�A*V�*D��,�5H�0'ᶴpW5Tu���.�J<�n�e��� '�L�$�][I���n���V����X����3d���(�q+a��艜�9��n�ne�6Hwi��H�+���p���̺��2qS����UB,�-.,�K�roar��c����YQ�����5ec^:�ɼ���zw�Ҷ��+)�R�Q]a�2���ೣ��٘�d�uN��R�:�Z��J4_n6��ik�6\g�rT���Al��B�̖�چ�S\��p�ux�e@J|�5�"���3Siq�*�/y�[�����x?��`�e��F2���m�L�1S#,R�6g�2�q���6���:��w|�	�\ב��X4!�,��� �A$����@` ���%�xw$����9@�a��5a�a�m�a�<Ȉ{�������_g	n+c`}E�����y�|�S��4���3���E*���28f� �0<g�bÛ�o�,÷�����h�`�Ï��A�9A�z��?��L����s�r�K�9}ǎ��ų�q��Q�;y_�9�����������N���3�}��Ӹt�8.p�kd�A_�½kp�y^���9�|��~{�}��u2AV�����y�A���<�w���0���F$Vb��cܸ|\�F����k'��Zl^������Mk���yc1g�@L�M=�л��*B��4��G9A�0Eى(�NB�����HT��b�оX4� ��}lۺ�wm�G;�`���a�:lټ[�lb%�~H@��V._�Y3�b�ԉ��٘?w���b�̩3~���//~���Σ��^�H̞��?���.���F����k6(��%�}���ǅ�wp��#|��{�X�	�9E�1o)�}�#����Ү�����M�q��8�-��A �*�t�z�max�+0�Y��* &��~�	g�JUz�_�|��<q�(y}g)�_�"��ևP(~�u����9��9!���JFa���
G��)�Q�4��c�_�JT��u&+&DHH2��:�d� ��r#�r��T*�.0,��čA��?���C��>S9B�����5���X�k�����.�{HR
�Q�o4�Kk�W�EH��ERF*�J
���mzN&���1ǡ��� �"D���T�f�}3�s��J�~��pp��JL (&��
�z���C�sX:��q�;��M��p�A�iW77���q�M���roB����7�%��Q��X�}���Ey(�넇��æ&�g���5Օ�0v,F�Ɇs%|<��`g���ɉI�GDx���Q��������twENA7Ĥ��+,�jX^�`޶PE+�^5�J\>����&J	"V��`V���.3�6���Ƅ�a,YfJ(2�;&#��X����	[��$0Dr�������j�3�e^��
Y��S S�ğ0�c�,D�<eBP 1��ÛU�F<�@�A�׬�1I��s�%�L�\�[V� ᳌�-S#��Y.ۋ�τ�j$CH�?�td�"�R_�A�߆�g'~�r.rnr�z�bQ�@�)�$ߞR�����^:�Q����	�ϝ�Nh�}&Pʲ�|':�\��s��/���\�@�_����?�ۏ�& 盭d"�ɡr�ٛ�2��F�L*�J��w*�|�a�s�7�:s��7(�ۥ��7�L�x���W::ye���x"U��^Y�Hu��:ɱ}s�I���7�~Ly���D�Ԏ��]�e��l߉���ƒ��y��5��c*qZ��"�;$�#��$Dw�߹�|���"�y��9Y�K�q�$�����`�W`X\�s����ᑄ��� 0lM��;	lJ*�o
�&o��r�p�r���|��z�7o��K��EXt�&A�W�������֬���o�o�����Ν�e����'q��A|�o}��ڡ҃{D�����t�6�ݾ��|���������ʅx�<l[�
�>\��6�������b�����G�@, �'�G�eX^�_���p��ĭ+_`��u8s|��,������>�Gw�������pl�zܹ�͟���bTcw4V�OU	�����Q[���幄�D$E)K���s�Z�����߅�{wb��X�t!f͞�iӧb���t��i�7�]�X����k�[����a���شa=�oߊ3g�`��-�>{.���"���c&�Dlrz���?=����u�0dAz�j|}���]�*���o��<�����߀��R��6�>��S�QX��8�Y�W�>܏��~j�����%H���_MBS��`��e�9�qb�X.MH����Ǯu�|݉@'0,�~y�f���׷��'�BF�W��p���"(�	�}� �W�EX% ,!��2S>R�p���|�z)?c�>��Wk ��?�����I���Y�K@X�a�3,0,�+@����zx�5�pm�BE��*S�H
�W2�FHZ"��W���l��D���#<|abn	Wg8�9���o���tD�.pvs&$z���N..&�GF�b�:�i
0����W��~C��	�~��E\L$�UH���&��j�b����KY~���U����P�2`��X@X�a//n�`������X*F�l7°���� ��r�V0�������@	2j�5L:v����,�loWgG%/7��'�`��&�-y�ai�K�`�y'�-<.�P>o�06=k�rY�W(Ig;��j=B*U�H�8-�K�F"RHg8S65��d$/�%<��7"����iL��Y,�S�1e����uB���/�Q���� �
����� c�����O�}o�Xu��:L��&Nt
��,�Jby�,�J<'c��\�**�����X��*چ�h�?�RVB��O�m��n�Ru*�yQLF��a�n�C�W��1�Gn�s��S���F�^2U>�S�<3�i#������ KM0�ZI�Sa\f�%�f�kp�Y.�N�\f�F�5!߆�M,3	z�AyT.삲��	Ǡ8r���)(N��%˂��̆e�y�m`.y�"�[���Ӓ�K�g�c+�����b�ΒPo�T}��F�\��M�Q��f"�2]�D�()���^�;j�k�Ƙ��Ae|O����kcTW�i�CTcE X³I��&�����$�p��������T �D`��K� إ���`��.`�]ö�a��0#wL�������`-�w���A���eZW�~�2�X����k���X�a#�<ׯ�R0|��]ܽ�t�������Q� ��?���Ϟ���/���ߨ�6Z�M���˸z�f>}DY��?��G�ġ�qd�N�6�flX���[?X�W��g�P�$�ŷX���^<��g�^�`��]�jf��O��R�a� �
��7����Ұ�%!�%�I'�+�?��;�ÅS{q�����ph��8yh>�xȫga����p�Tl}�,��3�`���T�Sa�����Y6f�ǔq�г��N`��wq��ػ{;V�^���Ƣo��(��BjFb������B���b��q�>s��;�cǿ�燏b�ǟ���u����1v�ُ�'b��[p��'8p����n��a��ۧؼg���ǜ���_�wW�@Ja�6aϑø��1�^��n5��j9��;�p}ǏG��)8y�1�� ����_:aGB{U�DH���8CLaV+4i��aB�į�1�H�S����[F��/%�5�x��V�阷��OT:����1���!�e\-̣���AWzˋ�[\�H����Rw��O�qS�#Њߢ ��'�7�3�"�n
J.�t8�0��vJ�=Q"-h�&֌Aрw��u,�*`⟣���S'1{��X*Nu��t�aX|�"���Î�a�mōC`X:�I�t��X;���Yٵ�a«X����D�-jR��B��%�Pn*����:�L��>�=.#VW�-��f����U����j�&� ��]�WP���:�����E%E��Z��|ߊK�Q��>}�`⤉���q����!��)>���WXA�._0AW�yQ+V�߸����}�K��GDX⣑�����4�FG� 7�i&x�0���P�)�I�R�����ظ�7aփ`쥬��N����ٗP�M8�S1�c#�i0�R�0!�����̴�����xa��h�vL��/)1^�fO�=p@?|��}��jF���WC���h�?��N@C�H����?�>2ܵĜ�3�Y͗S|kE�5�P�74�E=5%�dc��s�I6�T'�d��D��|/�8-�.;cɗ��ZM)�(��L�(�Tن�ܦe��:��b�ƦS{Wz���<�ņ�=�M��^FFS_N9ǔ5�����kTi��C1%6N���Mr�ƫA2��Q�E�ˈ&�#5V�z)Ox>��=��dHـ�O�����:���e,���C�}���gcYR�����L�^tW�y՟�-�2[��Ȏ��ω�fˆn�r΋_�.�@�����k��d�L]8���)#�I_���S9̼y}޼.7BP*�;� �a���O��o<"�����x�g�=$N~Ip	H�W�A�pʀ3��%$���*�K�S��F��ΒJ��r��H^�c��$f�3�Ǚ���o���%�5"�GR}�.qÑ���UȎ�-���k/�]�z�Le��V,�m���9�7|�5���FF� 0K'Eiu$��5M�p;�h�����/_�n� 6.�����>���&�$�'|W�O°7[`�Y��FG`xax�RG�c�0tHN�%+i�a���a�R:�8�T���W �zݶM&<M��]�S�`�$i �~���j��a�4>��J8gV �� �_�
�V��o����_��w�w�����
�<x�`��Ç
�����[�ek~���`%��K�����{x��-�O���Gw���s��^�������
�/�>L���8�@�ԑ}8st�6}x�Zw��i|s�"�= �>��?�%���KT��o��w7U(5��o�H��OE�&��K�`n/0���/���_~��g�c��%<���͵��l�j��0{6.Čq}0np7��W�1M՘<�S�Wc�2LZ�Yc��c�$\>�����Gx��zwc��wQ[��5X�t>�<�;����<ħf��b�UX�Z./��ʮ�ѭGo��8KV���k�c��X��l۱�;������<W�c랃��.A��Y�K�~�׾{���������cGq��p�.�� �(3W.Ɖ��`�j4M��g��>~ĕbυ���*�&�;x�݆" ��Y��8���&�G`����yY.�	�R�@��-�`��4� Ó�o[� \:�p<
>%#��p���5��l�[� ?.��
�1'��D�����%��@�>B�Tb��b+z�%�\^�Y�O8�p�#�Y8WÓ��+'w�Ra$T�F��H�����0����b�%�'T*e�UJ`����Z/�x"#We5r	�U��eJ>Y���rb���A7$��]���������&�>+��=É��'0�Y�=�N�ߛ�_f/��@-���p4[��ǉ0���M��WB�³���#f��}'�k�A���)N�8�`������q��a̞=[�nťK�Ta%�v�?��t\�"7��6H X��Ph���e_�?AX���+�ł����d��D�Ñ�����x�x�!%!9���� N�#������,.S�Ӆ#--���� {�s��GXH��C$1��2����F�"�s[�Ef*��ĚlogsS38;:�X����^<|��?y�Ǐ�O�^���@Ff:6nZ�G����+����=ؽ{>��#�ݻ�N���S��}����ݞM느�z�4j���5�?o`��r��|�� �����-˲8�M�P��������=�iv�f�e5*9�_$n�|_�s	պrz�%�E��"��j�-��+���v����F�d��sF_8Q�J�p���D��Yl���i�Y}��u��W���L����<\�y��}T��M��zc� &n�i�1!b9�j$g�΄q'JRg��3Nlt�u(O$��$�G+��L����2���a�H�0�F����T���t�]�|�#��s���q���m�eK�S���e��d�c8�P�'�H��2��Qmᕌ�����7�}ǡϨ)ȯ��OT��JQ�8=�&��v0���"���{�Bà��5l*'"���9� �y��R¶D��"��W)��,�����Y��Q��Z�d%Ú��[��� ���QU�d��"���S��>Xư>�y�ƭyl[�"}�6���X���W)���^����
�;��<�0�1��C`�B�%�{��s`P�r^`����2u��dԹ��@ V��%�@�1I��)8M%�R&��X��ؿ����s6I%��)���D�H�.���;�Z��a���1�
Y=�cβeX�f�m�h�ᛸI �s��{����4��o��?~��Ϟ=k���Q�H$���=�^�E:?%?������0�Sb~x�:�ߺ�;�.����w�
�v��95��ͯT(��߇w���7ו�XxrO�㻪S��?0_�8��Yv�Y:�H�?ݠ��^�)#{`d�
�U�a}�1�wF�ɣ21�_6f�?Z;	WNn�ݯ?Ǖ���Oq��Q|�w�*�����$&&!+���� �{�����($ ���x�D�7<����c��#�����|�$�sY&�b�G(J��a����v����6�=�wWo����4qVnۇ�'.`֚Mȫ�b����C�I��s�T���)���N�Æ����O1k�'��;�)Մ�����ʱ(��R�aX��°/aطd4׍�O�pV�`��KY`�5�;!�X}�L������� ,�%f�1Kl`WVTn���������]:�� ��+��JG`҉yz��#�xay�����I�﵏����Y�'�0���=R����¾ٽ�a�>��@J�����:�����*,˕U����Vo�DL9a8�A\"Z$�7��+�Q��|8&��n V��˖�Ųū���b���ݫ7�.YF��=0o�|�:u'O��ˑ��w�K:�	��|��A؏�'�+i�����2\��EHko<�s3�qy|t����!LSQ�����4dD##��&%& #=U�%6��t�sZJ2�b�����xd���3������Û�K2a�����	°��9�,,<�v-�9��x�����Ɇ�����7x�`���j̜3/Ĳ�1l��9Ӧ��	��e�x*�!$�����w.χ#=�u˘��������F8��4e,�(.��� ��7�C$�����{ԅ�il9��PjQU�F*�]��`�y�x�Aa"��U0�T���̏��F�9�7��� ��I�/�H��"��Bxu�6]"�`J���i�L>}+��w[��fh�Ǎ].D�'�W�G𚌦�O��Y���DrlM-.�W�J��5��&���a�C��T��rb��9��
A�,���T>���R9��0��H&>ٰ.�%ϊ�&.�~�x�.�=G��;8y�1�����C@\2�zc�'_���{�p�!,X�����W���;���Cl�wg�>(��c`���B�E��&<V�ҹ���+���
2;�F��O\�tp��
*j�V>����պA�h�����x�KБ���Qg�p��7�C$nq1!�VY���$�qSK�{��t�#�ʐ�up��!��7�0�-�a�L�zl�2X���o�7�p���0���ɭa؆0l���1�Y0[`������M_3���;�w�� ��W�鷭aXY��Q����m%�a���?�|�?�|D��>��Z�)W]*Dڟ�?=U!��uI�a�L�%X����g�O��+��޿��6������?�p�<�
��zO�� ���]1��T��A=�0�g������՘�9c���0�5a��W���{������'رqr��ѹ�[���~���[x��������5�ٺ���h����x�����#��p���O|"a����t񋅃W܃���,��$�+*��+�CJyo�U�Eje?$�5"��7�� �v2�#��	1E}��)UC]Ԉ�����=�E}[.�qG �-�����o@B��
�B
��/wB��%46 ��a��0l�1��G�G�3l{��<�Z}���C4�p
�ER�q�CV�a�������",���}P4`��Z�؊Q�ɮj�9_	�C�(�I2��N�t�H�S��R��@il�
��C\$<���AX��[s��N��`�[�a�+#��Z�a�W��}x=ٍ
��ˇ)7�����	]N��m@h6�J�_d�Ҋ����ə	��������VV6���CBBrsٸ�z''xxx�Qݴ8���g����ϛ"H
{{����i���$'�tS��8>&��	��d���J"�f�3RYY�f+��⬌te)�cz{�ßy�9d��%BF�	FH` B�����j��a�i �O�����-�ڿ�N�'�' !6NY�MLLЙ�Щ#��N��ln
'wW�����0�����-L-�����T���%4�!���|BQK�9�4�t)LX��,�,��?�H*p]�F
!P���;����v�yT.�	�1H�eY��� ������d�@!�K�|%�MuPǖ�*��|(YL;n>����y�w���=��W�I Iu�i����wrӥ`�p/d���u$�������Lܖ����+�{I0R�I�^ϩS ��N�2�}�w���p<]e���o��_�A�v|�s��Gg�d/��|�s��iNu��kaS�X�}pMC�TX�砋{������q���O��'΢�G��q@FQW:q	��;�}~�vÕ�/p��3���2�o=�	S�CL21nQh��N�I���tVJC'�>�\�y�;���T�55ð<��!�rO��U˼��%mO�;֎�����}k�$�l�����Q��!_�R���ڝ����[��l���ٰ���W�H���°��bQV0����é��d�:�@8��;� ��E2�a���pH��k�!7a���o>�k�n��[����៾��
`_>1 g@���_<�G�K&�Z_�_r^�����60���,���(q�_�����yq��7����˔[ģ;*���/0��P��5_c֗����oV���X�n?��������p��N����\�O�,����0�A¨e�_m&a8����1�w&��ܱ5غr,.Y�{W>�U���Op��>�{o	+�HU��Yڡ���[��]��{+Ott��l=��"S`�P�yG�52Ρ�p
I�cp2���D��32�1�O,�oB1�S��Gy'��7��S�1�M�-����"�g�Fp^e�L���|�+��*��3�A���C@~�ÙGb�x�U�Gp�H�F(8�TFV��Y��kaX�.�H��y�K�G �	d~~ţ�=�qu0���[�6��T�ה�V�VdD�� v�%+a�Gr��\��zx�'O³L��W1��-DR�8�\�Dx���g�Cd��Q9�}f ��X�]X`�Ru�[qw v��PrI�"���3�����bn`��"��G��$�wF/��nߝ0\�+a�
.q5꼛�/�)P��aʿف����c���L�I�ALa/����#8	��apv�z����Dhp"£���'Gx{����S�����Z���h2�b�r)m�M:�7	�*�'�a8��A��Р �pWG�F�!:"1��H��F!8�����B���������H�&���	�qH��_���
n�O8"�g�S��' N�v'x�� ��DH�S�$���R���/^�����-��o����a�!
���R�S`gg{{{�0����#)5�Q�
	A8�����7\=���������!�d�2���@%����c�X�D�Q5Lk�%XO�%Va�DGY�Ѩ�RR�kYe��)I|!�ӯ%e�,��I���D�(�
i1̹܂歷Z'!�� 1����S��Q���qi.����-����y�y�H	W�}E�	��f��s�R5�ù<L���T�A�L��Xj;�����i-ܖ&��;�)k���.j��n�{������"R�ˮQ���4Ȓ秩RI�W�����e"�N_"��Y�V�c&�� 5o�X��c�y�y�´��}��}�$�[� 	u��lpX�qcIY��aM��zS��_ٰ�v6�Y��9���\|��Q\}�#�-y�������iX��#\����>ű37�e�1L��e5������0��e��	��l*��|�)�;�﹔w�^��7囫$���{/������}TGR��'�_ZGL�;ʢn�I��5��6��̹�Ȍ�a�}�	>�΄_�4���i���#�/<��Q�-�,�V�Y1�}K{f�NN���|��Ў�u$��mx^����EXN@�`�3��U��H��a�0�b���a8��e�6�i����"� �K	��0|�0|�����j�( ��t�$�>"nw��xN ��	�ʭ����Xpj��i��-��ͮ���C(�ɫY�:�b~��=}�^��:��/����#X�pNނ�_ħ-���������-àt����Eސ���٘:�s�Tc݂!8�g.�ډs'v�����t�V��r1��Ю�):�;X{��c �����	��B����;�@������d�&��P��"��xĔ(�ǖ�-��	��J�"�v'��GJ�XB�D$�"	.��]1Z�lx�h��(���CT�$DTck�"�v!k""�&p��-�v�䘚1���P�D`����誩�������+����.�BMV�aX�%���a�aX�h�A��d,<s�	�Z�>����%���ގ��¦y�#Kx3VjZ$CLSp��',�a�8W�w�G,C��e1�$<K�9�.�7�U������r����Ab���&�x	�pI",�2��	���s Fm	��􆩄�z�Z����ؒ�0L6�� �p��i܇0lp�v�u�'W�/� =�`��y�4q6&O����`�ԙ1l$�[�S�LCCC/�;k�~��[�c��Y���C���&#��(n*��q�aX�O6��f�a�t���paA���!��FHuQ�+���i�\�˴(>:���'�J�Z/´?�٠�!HKx67'�<��'|=��!�%\�H�6?ه����wBL��a�̧Y��	n^p�s���~��������j�q��l��C��Q����p,Z�_�?����aʴi�9{��ok�n��5�ڭ���Ct�;�]�w�+�������o�6��78�?<3�)�J�H�L�e�z�tٯ/���<��}�K�q����}ب��zQ=�����j[��>|��@�C��	�4M▣Ip��z�A��)?��k�����jj%Y��k�"tx�6*��u"|�<��Xm}�=3���<r�|�1��U�ևjT�K��F��4�9����Fubl�ީхp]�hwMi�L��%�I�����G�H���\�\u�L��2�;��Z_	���)�eWl9�r��Q�ʆ�Ѕ`�J(ug��ZǐLe̙�`5���#�́��܂����f��ٯ1k�*�ݴ�?��_\��_b��0l�Bd��3z�!�,Cs��P�x1��gq�T��0g���Om�W[:���s�&���!C�Rgn�d��|K:sJ�L�sgK'��iӎu�]|%�����|��?�wS,��NB:���.�+:	Gt�;5��C�U�=a�S+�s�n����0, �*Pl�~�`�@���j�O�mn��+w��Ǵn�'F0��}�7߸�_���w�0,k�Vb�v�u`�g�����n]=���F������O��pMkB���J�����I�0gT%揫�����8sd=��Oݎ�7a��9��;���������#����#�;�(�/� ��s�,����8*P�L��O:�K,�"�o�&��ɨga/�Ew��%؎B\�q� �	���o�8�cF �No�c�cX:~E#����E#UV9A%#�_8�%�\6B�U=�%�(I	��S��	���0����t�eX�dV�2�����h4<r��:�[�l���V���A$�d(2{�@R�	��+1��%�Cz~�����[b����	(��u�[�Da�Io�:�#,�Ȗ�� O|�����k�@�7+s͵@�t@��r�!���]	���ܛA���b�"�V�T��ZM`8��X�{�����]�3�t��+0,�a9_��@l�1��Ե��}S�b�-�O\>���������g'q��|y�,>ٳ+����W�)�a۶�{�>��8~�z��E������u�<�|x������hd$'"%>>�
~3S�������B�e+@N��ABt�!�jYLD(����� ?�x�",؟��E�uV���X�؈N�1�`�L@�`�ߛ�����#ḽ�����"�:�����3���$����m�mx��1�u��n��O���?�����|��il�q���EJQo��!�^� ¦N%��i��{e�L-ז�|r�+�� �,B���a���w� �Ro�`����`�c}Z�$�D*��Dh���R��T��Eu�$���L�O���;�ǝ��ؓ��DBlbnÔrK ���(WIY�:S��"��@I�& !F"Y$�.�XN��?�˕��۔dZ�m�r{����`��c)��z�59�qM��\iP'$�J_�u����j�h�$ˤ�\�$��.��<#9���r�qO:��h�}=S��(�p�İΣr`��,��'��=V4k�<����3�n90uE�q3���;h9��a� K/�l�c_^"�Ĳu����Y�Z�#&/����c�ᯰl�~�fT��[,���{�6<����r���n)l#+X�U��嶄/��׉Z"t�*�������wZ$	��h-��qY�nPb��DI�9�@�ˊyXq_%eu��|d���pg�H�q",��!b���J`Q�F�8��gX,��&�[�ŗ[���gK�֖a��f�&iK4	�$�G�Pp*n�@l�n�O�UN!����Z��A[°a�-�[����`���;���}�%���������`X X����`�Un�]I~���c~I��΍�X0g>ݳ_�ڍ�;W`���6�{3�!3"@�=��b��:,�JM����g{���-8urA`V�Y���lt�v��[0lS���L���}@��-o�e���}`Q���p#�@�Jb�F�UKdTU1ф^	s�7 U���k:"�!�];1ݧ �� [9��\^3AU�M��קt$�MDD�)�2��x4Av4B���T1��'�-�h�O'PO��a�>�b�+�Xb	 ���q�)����w�x��+��8>\>�J�!�$,>���]�v��ʕ2��,V`���r\.a�!�Q<U�#�d0�JY1ZY�K�]N0�Dh� d����nc��^�(��XB���D�� ��.I2O@��PVa�a/Ð�
�	�y��e8�z�g�yzg�&�Nfa��ᥬ�jTh5c���F�sM"��i��^Ò�uE��U|aJ:��g�BHn?D����ٛ�t ԬC<�i@Tq�*����'���*�zn0}��Ca~�,�%%e7n6n܌}��c�����pttT~�� Z��n��A5t���V�ᨰ�b��JKFAN�]�Ḩp��9���V��	�b	��D����i�NOFbl��]�u��ȋ����DuuLC4���n�Ѐ@��	���@°7a؞@`Mw	gG'<>\�׭è����%�
е���Y�o�Q�G���S3������ZT��GzQxG��.0�A��ݓ�,�*�{��"P��r��r�s�Z��"�^:xIg��U�ۘ�'t�m�Ԋ��2Me�	�G���Zd��;�V��T$#��yʊ�e�O���,�_��K�Y�E �,��� �U
��2��)�VA��Z�*o\$�TT"���DP��y��i�UBS1��l.��梈2h1~K���r��}h�����%�� n��2��M̂���a��SE�n�Ħ���#���6�$&�\8�x��~��о���*����`�@��a*����磓O6:zg��O:���dt�N��W*��2��G����fA��	k�8tv��YKp����=|4޶�E{W8x`��8|�������)�'�ptq�AdVVnۏ�.�Ev�����ήa0q�$xG��{4:x�Q	�������h��Yh睭��'GIK�S1�;#�����Y�?�:���)�~��}�;��0��&�.V~��/�	�_X|�9-���*�5	��	paCĕ�9�mxa��0\��A�!���j-�#Xg�q�0��t��,L��:k��4V@���g���pj�k0lJn��`�κ'�V�p&ax��eX�v�l��j�&��{������G�ZG8M�Gk�@�.���������ʲu�1��ƻ�6UWD�̜������,�R�)f�e�L�2�l�Leff&YlKX�����?�>�)Yv�U�}o��1�CF����W,�@9����/�<0l��o�_�'�G0l��RP�.�/����O�K�ᦫ��+O݁�؊._�-��cxj=��WaA%RK�Tc��l^h��uLõ��mW/���^�瞾�?��>q3���JԵ�Èu" 1��j���l�N��ř|a�����(>�q!l��ٲiTz�Rd�-CV�rS�ͨk��V#K�/�W �g��7b	�Tv�&��`l0J�s�R6{�ZNכ��~'a7�k!��9ur���qN�N��*�� �EHUМ���n v�`�O�ѡ��;���m���5Hm[�Ć�-�ߜ~�j��ʲL&�.AӼ�����n�a����B0,K��)�v.R�g���k��UƇ��&6\�H�����V±`�{�e����@����Z,�Z��l�H�<�	���R��2��ѯ��	�e����e(X�k�!%����50ÁY���Q"�nU�#��v�V3�����TtCA{9`�:�k�j,`W��+ϰ��us�.�X�b°,z�>ſ-��-�-�Dz� 2���]�������@Bb*�����hClLBB�O�u�����d�X#&&�����
^h*Vn_ G�MUe����T ���'�$��B�q� w�5ȭ�(A�	f0��O�q�lM�9N���Y�	��]�
��r�}�����墈P,0������QUV��t�N�"!�
Y��Ga���N����_��̌L���7�����!�?L�8��q���0�9n�����:������m�"L:덏��=�O�#_<]�r�a5�D������I����Hv� 5%\Q�! H��N��[w�x_���~�Z���l�� V��j�j���_��'��_j#�-T+�S�,�5mG��P�$�;��LEP�̔��6����wt��Y�*pn9	�����V�2����T2��H����%U���g;O��T�$����jrK��K�x,�=���7fm=�%_ʏ�$s������;Uu9U<SZ/�T����R|%7+��zL$hN$�NL��m+����0\[!���0!�>����*�]�����f#0.+6_�W>܍E��a���8G�0c�rË�lB�#��,L��q�шI/�ҳ/����Ƽ����l��N�Ee����K ��=y%�	�^�Z�z��7�-ƯD��h��οG���SRU�����U���<"/}�?ki�;xs<?�q���� ��y�8N�3y�3x�3%�y*��+�W��S&|Q*�����n�sM1��R��<�*��aPTzZ�=���*�p9a��/����40��] �
��0|���aا�0\i��o�
n�	��qf^/B��!�}cl�������p�6�!��Ovb��]���=�l�޿��9vǎ�ǱC��������έ�	�#"�Z0|�0�`9��V�ܩa��������t&���Ob+�΂a�x��p�Ekp�9K�ؽ��q�V��[�b��V�a�t�����e�d�T\�e6n�x&n�l.n�z)�}3}�J<��x��q�-ע�k
c]�M�ccS�3ٸ�Kz?�1c*Ns�rT��\%���$>ж�%�7.Ej�28���ռ�P���@��(�CZ���v�E:�V.�ڌ�MFi���
��6�\?V�>B%�ۻ7 �k��z���R	�Bh*�3Uj��^|�.J ��ã�%8ոD���hѹ�?��.N�	�M�9�^���� ��Ӕ(��<�i��^�ꡳM�4U�	� H�*g�T+cD�L㋨��|rߊ?�~�9H�$vp��R3���m'��l�Z��<-����G-����˵�ñ��n��FWF(.�GB��I��iߙ��e(���JU4��\�Nو�J�����x`�y%a�-aX�*�	�Gs��	��\7
�Z°�re��=p@��jɔ�8�@�ټ�X�C2�c����rI7?��eT ���խ�-�Fqi���(-� ܦ�l--����FVV*++�������+v*�Dj�(���к�D�[jJ22ӝ(*�5�ooYqj+K	���b+�����r���2��.��A�s���v�!�����վYi*�a7n�b��Ƃe�^��Bp]N.+,��\_���l��:�߰�]�4�"  'Lĸ3�D{{;���zܶmV��`.9	Q��s����y睇��>ӆ���Ԍ��)h��Eck�f��wҊ��]�$L�
{�l��2�B������<��J��U;�|ܔf-ϒ��T�h���i'��-��gh�i=;��)v��<���z� )"��9�T�)�畊�L�o$��&��1��|���\��(���Lj�E�� 6��vd.a"��Y|�3�id�D$"r&#4��=&()$S�mBL������0�k��>D��7[�`��2Ⲭp*r�O�K�v�T��8Q#���-)�,���TH�:n�H���Y��T'0��-�k�r�Z���,K�gY�<��/��U)N�N爂$4UYnc	w �g@8�!{Kc�<�d#��%n.�OJ6�s��XFH��_\9�JFP���`�������һ;�����9�!1�X��<��^�Wo�9�_��V��xxG%`�����Kocڒ�<g:&E��R ����t��`� �ls%|Sj�4�l)��t����K�D�JiS�޽ݒaKM&)3�OhR����M��M�_ ���Ϟ}Ef���%���`̛��`��1�È�Z�pBbH�����	n�R�L�3^5� °�`�K�U�(�sçF=a�>q
�m�}�3t*����#�pa�ڂ�3پ��@٪!��_�����10|�m�፷�;��@��_;�����"��S��_~��ǔ�̲��(����)�,y2I�4���}����u�y����x��?���/����ykg�tj�'�`�d�g/��%�f��g�ƍ/�͗��-W.��W/�m7n���\����<u+�~�N�L�	�h|��9���|�-$��%Q�����$/!/%/#/'/#/'� �$�6ʔ����u�A�0�5�P��K�Ҩ�a8U@�0�m'�0�>S{(M�cd��=�/�a�;UU��ܾp:��8��k�\0���¡�����̩�q!�fnA�tB-!W��²� ���eV@�|��:��c�e�&P
ZC�[Mg�D`M֋Y�KpDA�24-�B0%�ӎTƇ<v�V���27�>�_�JoK��\��'��a[�c.����pt��%��C�B����0,0��p%�=��j�_;�^<�.0�YVc�UK��m�XU����h�R�fu(��<���ms��!�eX�w<��y�I�vǽ�����s/⺭7���4���w>�n�j�n�ٳ��w/f̘���4$&&�N�tU�͸I�a�U�d XnJY&�paA��\QV�J���%�(�J	əY��r
�塙�+˯�*,X��r�("T��+ؕۄÖh`Y>��O�,�d�s}u�2WJ�DEq1�Y���N<��4�0� �@�DǠ���>���ۋ]�w��_�����ю��:ܾ�v9|;?݁��x��}�~�Y���{�p�n|��}�],�t*z�!�a:R�*H-��Xg��T�2~�+���6�2���?Rz�
�q��m�QZ���\�</��l�����ִ�(]j^`�Ӝ���0.0.Ee�e�.�yp5͂���_���i=�����x��i�d���d��Lg[��v3�q9׭���ls5����l�橴�%��/�g��ܿ� ��f ���������"`�dQ���~a���G��wK���pJ�R*��
+n�@�q�R9IYrm!i��a�H��	C���ki_�m��{��:FE�T�� ��n��&�f|e�Lm"7��I��pA8��20�K�O��\��P ��4�`sʛq���㮇�Ô�K�Wֈ��a�������5�s�����p�Ȯ�GU� ���^����	�6xE�"ĖG�Ƥ��Kh/���� �_Ja��a�)W�|]MnY��%��wڨ|�%��%oB�Xy	z3Bf;ᙃ�t��[����Y�_	�`K�z-s ��e�)Ǽ*�!�$Nn0U�|���c	������5�z��/�WM(����P,��?�ǝ��Rq*��[��`ؿf�}.� �.���j�p5�'��u����Ç	�p��0u�s�o8���[0lItW	�-�1r�N����{�`k��ĖLyf������}�O�7_�箟�+/^�k/_��Z��VNô�2Ln-�����)ú�n��z*.�07^��_��J[W���7`۶p�W���n���<��)�1>8��uOqðR��K.�E^J^�6�M+؉	����d�ƽ�LeH�a���	���t«�F��9v��rð�~�!�-;!ԣT������p�)�s0�ڹ6Bp��":���H�g���붭BT�,�*m�R-Yi����e�/C��eh�{�^6>r�P��r�%��_X�2��}�(�[C��E��Z�1a8e6,��0o3jfmd�:���7�c�&( �H��c`��q�a�P�67�*�J��`���kɼ^r�tc.�I��+0<�9?ü��Re���XE<TvY>Ų.�dtDn����5
T40,����u<����O�Vn�5w<������~�����[��[���g���_�;�Ô���_�L�{˗/EVV�)j!�ML�7��r�f����L�b�U�"���%����C�XU�r3���Bvz*�S���Ǻ� 9��\�.B����!�`ƕ�\�{,��W˕���c��~�Vf�Z�pmE��[��D]e;�T�D' �;���+�,㯿����;�`�x��UhjiFss3n��z|���x��W��+���e�������W]�˯�[~�.ބ�V�py/����Uol��
K�UX~��12��i )�M�,Ŕ<ǫ���	�*���s��TW�|n���ThJ�_R��D�ȭ��Rh����:8��=vSJ%��i�a��3����nh.�9�9Л�wo�LCsy�*�4fY=P�0M��L�`�(-Y�qe�Q�ބ�&X.�w��w� �aY-P�`�d�����X{	�9A���Q����`*�X�[��ZG�a4��L˪h-[ ,"LK:����'^����Xޛ�1���h�Q�;��I΁O<�4�~1�"���?:�B������9������#x��ݸ�gq��w��s
�������� ~�u<��x��p�S/ax�yH�)�i�q��r H.�q����x/~I��M.s[��5�װ=r�Ӓ���$ ����J�f�,#���c�%e��0��J�4V����i�?wY�C�5���E% �'f��t������_�a��գ0\���G-����;�j����g=!�#��o����B��B��<��w�ق�i10<�D��?��:vG�|A&�7������[nV`{`ؚ���p�,K�( �3?�Q+��-�~��>}���\|��x�f<r��x���x����ݿ�]7��ۯ;wݸ���<y����sq��pߍ�pύg��6���M7^�۶]����=��L[���c��_L��ÓÉ����H&��n(v6�$�"���Ԧ�gk��:,L�\O�`8��0������a����>,�-��Q u<���X	J-����3<�zc��	ֵS�Im��|F��pp@�JNmY������؀���c����Qг�×�W�c�UX.�a�l�	Ǚ-����$�
����d�H�����nD���0���BӼ-p4���b����;g°�,��)�5�`���I���kY�8��˺�Di��k��,s^�r�n0�S2���y��&�T`f���u?bm�g�-2��s�#�e�q���4���J!V�j���� !��Wڃ����VD�#���i��+*GYy5�/�	�(..EFz�����*̝;^t!��ZL��x�iff:rr�,+pJ2������g`�fK",ˍB��-�	�#E�[�(-V:�4��&Ù�@M�4�-���W@�eңi�#�uB��Y���X�q�^�	��r���e�yf���Dq^R⸜�ֆz���>xN�w���v�����������o~���ٳ0e��'<������b��I���FiQ�)���֎j�\-�iH��#(*1�|�gU

&% ��$�9��8��ϫҙɍF�S�0��cMLm�Z,b�3���(�'�vv�n���\���hƙ<��ϰ�ڶӉK�%�~��ןak4�ȧ�L{ƥ�c����[j�r3׷p;�ԙ)-<���k����*Q�-<g3�Z���ө3�wۚxl��&�\�>3��DPM��c�7(8�`ۡ�r���a�˿/�c��'�@'���U�F���g�U;E ���O�lC�ӛ�gD@���ޟ�ey�+D�wK0>	��O�a��F�4��b�;��+`��V`�G�2����j�U�`�p@L6�	�1�|x�$�?"�M�ظ�Jܰ�!�_�~(��	��#֕���v,9�\\�A�9WnE������c\H��������,�>1�\·b!���Xߤ2Bq�b��j�����S��a�?���Oȏ��g>V?b��]��'�r�8Q��ٗߧ��i�Ձ�/��s��I('k�W;������0|k�[��0<
����6~�gpP��n��b?U;��i��U0���}M0V^a+���Xb�p+����(�kZ7�=�unM�a��:��Ζ�:�)�?Y�X�=d��N���~�/�'���;���	��8>��*�?�	���x�ǽϿ�C�����	<�ǫ����;.��w\����l���x	n��rܲm+���C���qA����A0|&a�7����a8d,7.3@,���Av6�"�6J#	�ݖQ�]�@�i�2��0L��\g�� �1 ��$V ��
�K�X���屛�ѷ.�ݶ�e�������lzΗGI͕v&�T>�g�s��M�������	|���58<��P��.1�&�aXe���I)��8�O����9��6|!l���`��ׁ��^���`8�̲k*6aWp��+)ϰ�anWv��JYg)°G�]6�a]Y�=0������kG|��M¦ ���?�ao����R�)��~�\�)k��3�E}����2AsJ'�gU����L���DX.;�,j���	A�\����0D�%c�D��'���aa���4����8q"�Џ�����2����i���c�����~H'�ْ��N.*p����O�=�FR|b���,`Yx5��EB.c����	�5�()0�r��T ,�
�G� �Y>�V��|��"$�������2l��0l߰����>>���?��?!08�.'���Ǐ���$"2A��GB\x�z�	�4~ƍ������i�1.0^Q.x��"$��Y-�-&X~�9��Tt���������ʸ2`��q�*V!���R��6��Ȏؔ &����󖲹��?�G��� ^�� 5���Gij�s�P�9?�ȏ�U�dIr,iޒo� |����7g2���^{��Li�ʞ��־F$g��{x�*�`M��2>���n��p�9d������B|�tk0��(3������O�ɒ�n0�r�584mTa�v"��QV��`����6#A�1����~��	�uF��y~����G`�!�@'�aOrð7a�W���$��'��0\B�GP�`� Q��O����OH��Fc�_�cR������/g�Drm��Mƿ����h�;���A�	�~��\��iU߄"�$�'�>b�dˇx��i�p a8�$ ��RGt �*�����ܞ�V� >� �0_���5�6��- T[0|&ۍ�8(f�~0�0\=��&q�-7�����ǹ�0����/�՗�L�5S
���8�^%���;�[��
! 6�<��1�0Z�Y`k��������ׄb�d��f��]�O�oǫx幻�����?n�Om3�o�� �l��z��|���c��!<��{_Ƴ�^��n� �z>��"�R�sە�㖫p��7\�[o�=�s��Wb>�	��\m��S�pB풟�a��Pܺ���aJ���y�$��%��P>i_���)AX��H��>q�vJ*�|��	�;	���! N&;�߻�KH�U�'��[:�D��j桨wJ�7"�y��S/7A�,�f�X��Ia&�Z���W,xac��i��o��ͧ��@ٔU�"xv-F!�'�
�����[�a�nV0�@T�	n�'P'ð�K�Wz��)+���)�sِvX0ܷ�=�F`8�vʧr ��D�'��`8��ǲ$O?53�69`M��h0VaU�S�L�6ᬝW�$���+�6>��-���r3f-߀���b�9`�aShchh:��[`488�ٳg��jjy2��
��AuK��,�muu�q%P@��gee�	��3������ނ��
��W+�wX��BR��_�G��dY�e	�k\c#�6����G\Q\`�	tuN�*+2�²�|�n V!suY)��4>�*Ǭjtr��@��~���!&6g���=���Eܺm�I�G �����+��#���G�m7߂λ �]|9.��
\��k��ҫ�|��h������j�����p��ͧTpc!R���|���/Dj��	r��36jYf�u��r]j��4/��9]�d*�yT����s�Sq�N\�b�6,E۷h*�~	��u�"3oi�[����H�uy�Ė�F	�˸~	��\��:>�Fֳ���Z�Hv�#��r�B�<���A@�4x�&�s@��b�l��U�2e�I���vC���M��w`.��Ƹ�zx9��6ᔰ$�
$��H� �G�:�Xq���6"����ŀ0�Ib�3�Ml��+��ri���:`|���J�F�5 M�2�ʢL�z�.��I�}�2)�Yh�ľ�>|���EXj0!��	���119^�\�p6�3ބ�PB�Wa���%L#38�Chb6�Se�؅�}c�nG|6҆�x�+:���>.�#c1):Ii<g���O '�������Ia�'��v���J�7�e	�D8�@�'����@�N>�����]��������A���"��|7"�aU�F`X���X�8��Ӡ��XH^d�I�V)��*�FA��+�NnN�B�F�(��0.�z�	0lR�m�����<��aX����J%$w<w��;���]������}���0���Vje黣Z/+��=���;�+YV޿.�o��ax����������G�e�=�	΂����8����^��x��mxU ����޳��W;q���ؿ�E���Y���,~�
v}�$��b\w�j�z��r�Y�fl��b�u�ո��kpa��nFk�,��ʿ�Y���V�.�����i�f"�`�(�9��?Ò�ã�YҺS�4�O�a�O�a�����R����[֘��~���y�u�a�6�����.@���ѳ�j�R60�[��,V5��\���۱�+�F݌s;!��f�U�"��f���	��P��ٱ�c��:2��ed��A ,�`X`;D0��J ,�oR�4��K�{$8��ǖ�;��G����S��60*_���gX�8<0,��$g�/�����U�
�lh	�r�h_rjfn�g�o X��h�H�K�0Vb�]���幝�P:��ku:�7གྷ�aϱ?᭏va����|�A|���x������o⣏>��l�Th�~0ҫ���+�#/?IɉHLJ0>�i�N��բ��°�'��
�@��Yqyi1���g�8�FIaa����:l
��߰�X������QAW�Z� 9A���1�����.�;��9AoUy��
��J���:Y�K�	�J�F��4͡ :'B����WU�:::������q�����0g�<T�T����w?��?�c��³�Ά��[o��w��o���{�=<��{8�ڻQ�O�����yH'�
v-�U��І@wT�ئ|9+m���"ce�6;���XJm�2���V�"�x�d*���D��-+ײ
�l�b�W#�i%��lߢ���p���F�2��uF���yɬ��q�_�(�ud�3�ф�H�B(�8�d�r'c|z���:�p;��j`8��{f�J�cbJ����T�wp�	�'W��Z�z˂��S�p����V0�W^e�	+����7�X�2�	8<G.��%�R�9n�U���I�`X ���(���`8�0e,��/�ϱ�-^S����]���\n�}��)_=�)�Q�Ap=|SG�>v�EbBR	�'bBb>&&�bA�+) Q@��^��	���2��Vb\�A�y�H-B����i���S�p;���$��7��D'���Q�8#<��i��O��6L�q~n�|�s	�yTUd���{�J,!��a�����Fa��*a@Xk �����k��/� ���X�GA�cm>kТ{�G���0�v����aI0��j'[��K�[?�&pΣS �ߣ�k����ɖ᠊�e?]#��"\x�V���'��_�3�+`�(�>@������[�ٯ����Q����؁O��aA�j�\Yn��z���v��W�`�s��	�c��1A�x�s}}x�2>�ò
�x��0lY�w�}u��_l�����	��î����w\�瞸	o�|/^x���ʣ������x��pd�K�|�ӄ���g/���W���������]��n��^�7\y6n���~㥸�?��m7���gD��o/��[�������M���GΚ��!B;��eF��G`X~�&��@�*vV��l����վi��v��#�u�I�<2�J�<�d�,�w�����7K�4ͤ;s�C�X?�T���O���zr�����^'�� ���Y6�R����OVĭP5M�z	u��?��\���HNc��PB(-����)\?�����Q'�0�Wc1�����j���P�<w���s���H�e-VYe.ǖ(�p��7���
�3lY�TLck�!N��!���븎�I�b7�"l�PH�`K��7�D#t���.�#��"�2ૼ�r{P
�ph^!��=YkY�e���Φ��zl��a|�e]�<s�N�'�$Y��yD�w���p5�KڑZ݅�W܈��r�ބ%+�↛n�ҥ+0y`�]z.��r̙=�_#���ڳg/�x�I�O�������h�*��[��Y(��@Ii)�J�QSS��Rp	r�3����*�`����$Ą#.*�o@՞��pS5N�_e���ײ�ʊ\h Y9k+�Tn�Z� 7'Ӊt��Lr�y"�E�`��.�br��eX~�.���J���|*�CB�珨�Hc�~��9h�����`�#,X�			(((��W_��|w�~��Y�v˭�2M��2=Cs��Ρ�w��+h3��+��V�B$��<�PF@����M�[J�>ss�w@�!���g��z�����j}����cuLB�lD��Y��x�����;�����Ϋ��?a<�0�B�e�ݼ�F�I �l\����r�H�wR���H�G�sY�Kx��>Q�j}�G�����7r�[��^� ��sR>��3���c����{
���\�J|��|�Q��U�ᴸJ��V�.IJ�  1 L�%�Hf�,��-�!'��8$�����pZ��� Le6��	HPN}2��2����j�9æ\�(��G0ۅ`���[Ve�'x�s{� ��W7!�~�$/����u��^�
�o%�?�Y� W-�S9�����TDb�`��;)�0L0�WbbL!�b�)��b{fD�6���G��AtZ9"��`�l\�!����E���y���H���T&�fRY�"����;��[�J,�=��ʌ�.!W� ���ȿW@�϶�ӱ�M��F�D���_&3q[�Gax�Mf
:���n ֱ�a>;a|���uK9�FPj�&�a=c��R�y`x,�@0�T�)������+�G�u��آ���`8�b�*�"�z*j�/�E�_�kn�e$��/��Ç� �`X ��ߎh�����a��c�	�V)f�@���~|�r��]B�7�ey�c�^���Z�<��AP���~�c���O����Gt� ��'#������{* >��}���Э�xn�X����>��;8~�]<�čx�����3w���O܇O�{�����]/ⳝ�b�O�~
����c��ơ�^��o?���w�|)n�zn��<����p�֋��+����GQ�T��3���Wj5_�V����TUqb'�=�C�c�S#��r#�W��!���<:	v����bGaxT�����K�5�[˞m?	�'C�	�O�^1�=�a��%g�Q:�0�L��̥����v.J6"�/��F��"��F2XJ���H��`G�ۺ��/A��-p��&0w#����)kB\�)Mܾ�"��s�N'��X�s�p,�?����Ă[c�U0\�t���Q7���l$q?�%�@0aZ��b�t�qm�
����aW�B�	���+�+��Β�`j�\��X�������s����\$�&�%�b�s4�5���Jk���eB�0e�P)�`v�~�н���y�J����'�����$�"00��M���������@�����!($����w6"*�0\L ���~�F�.ׇL
󳑝�2����c�l���������+,��	\�KX��J����l,���
l=�^���Er|$Ry���:�0l�p]u�9��4d�6��`�B��н��߰��7��_��T�KNNF$�X�G��������i�����?�'������?������ x���/� �뙓0�/���L�F�����r�z�6��)(R6�)�;L'��1֍�� �07ɡ��3?����~��dt��*�p����!)@.��'Us�*���>����&��,_�w���-kEE4�Ex�j���V"��G�l�<
#܆~�%AD���j��c�B��i��#��#$�2�ѵü'.�͆WF��a�ru�he�H��G�� �t:b�N����Q�ͼ�yy`X��S�_eh0�|��Z�"�܂0*�pNH%�~C2����\��L*�a� X��L�iQDp^��G|�����p�`�o+��PF���|3	ZT��9����}�|�~�)K̠��+����n$��%���8�{�]� >OR���LC\F�������Iyf�����pZ�ޜ�K��p&�L��!(9��������t�f��Rpzp&D�c��<^Y"�	��/^a���sܖa)߀�G:&(������� ��R0�8�)(�#��?��P�@����}3+�P��
v������>a2S�/c������h �g�� �=�ߟֿA���_!��`�܂�Z���7܀k�K���o�>f�I��:v_?�������,��a+@���]8�9����8�����)��+���k�8X���|�~G�ߓt�<*�[�$�v�H����AB�����qd��8���8���}����3������+�߉;n�O?~^|�������ػ�}����ᷰϛ8��[8��;�����*>|���ړx��g��]7⎛��]�lŝ7oŽ�n�wo�y�
9�l�J����#m5\~i�;{J )�e�+�cJ/�ã�V�*�"�r[�
��O{2��������܃[.j,+p*e�R:,���d�ag�`X�����rr�W�,�`��F�V�ήt��ĳ3p��CÌ-h�s���d�2�UX�I@.�[�°��*�ti=�����&�Ti�a���`����xY��P3��JB|�:�Α�h���{���a�0x`X5�Sj�Nk60���Qؿj���P4��p=d`X`��l_l�U�9�f��"k/%�be����$s ���;��!��\~a����"���qN+����Ϯ�r��Nv!>)�q�HHLF��	{��T���M@dD�	��D@P �SRPP\���B8�N̜ͭ�`XnVJ�D�fg"Ŗ����]��R[��nR�)װ,Þ`9Y�U,C�^Y��*����l\(�O,7A���Yn�g�����GNw$q��fGn��ǥ�kɪ�c冑N �9V��3�8&�Fyy9T`���j�R�{kj�������1�ѱ��I@F^12
*�^\[~��j����01���'�S=[S����]��ԛ�M%3B���+���T~X�����������ʙ��� JA��&E��*^^����~$r`�$f�%�lY��f�iax�)`x�����ZJ���u��kY���Z±�����an��]�(��`8�y9�"�h�������ռ����3���1EG|�;9 ��g#hQ�5����
���[��a+(.��F�
#��g5#:����s����8��BZ��
���}��
����(��*	�ռ���@0�E����Cā�{�]WN[���a^˂a�UB�fTl$<g���G(����W�o#tRd�u"�Y�AU!���L�E@R6�9�
H�A�� �b�k�9�rS��F�~��s�OE����+���!.����\_�u��pFTZ�x�@��?���3�nCl�ܧ���Z�R��+Z%�-yǤ�Z���%o][���Q@"�c��|T��8����sw�M�အ�@+������e�%غ�s0l��H���`Xn ���m.|vTF[0,_{=�Ջ���5�U�n��#��Dh�S�.@0L�O�X�$����0TFVb�]5h`�қnĵ�n5E7�|�]�޹{w���;��"��,�_	�Qq��a���0���A|ux?��b/��`�G��?��&���>���%��d�[�G>�hD����9Q��>!K�eAkE���e!�X�->N>v�ޓ@�]���;��&�l�_��ݎ/>{{w��ge~�^���cx������c���|�N����>|�����ط�C~��c�����'����ųO=�Gz�=��x�1<���x�����K�R�Bpj@BI;�F��'d&s(k��sŇ<�|�O���,�M+�ڼjD?�a��j=:����&&�&S�_�=���?��H��x°@8<WV��(�[�\�p;�ȼ~D�ѐ%�`2��O8;��Ε�+�l4�a���%��J	y�H����y�v��y��)?�A�F��V6��Fa���*�5A8��eY�sz�"�%��� �ab�*�!�."���<���ռ �k�?pHN7au6��4/DP��w#�k��+龬ry��^Cr;��ҫr̚W��`Y��C�de�б�^]�X�	��*᨟k��yW�|8�����K�9h��u�]�+n��\u.�r+n��V�y�=ظ�,l�z=.��R̟�K�,��߅�~W]{&"-#���'�pvn.ʫ*Q\Z�q%?a���ٙi��JCQAr8��*EEi>��5��gX��,*�,W�J��,w	�W:6[B2���B�Ǌ,��_8élN�.{"l���h�&Śtn:�rKiv�)͛�뼎10��_�������8��z�޽x��1}�t�N.##���s���w�Ý�߁[n��<�^|�u<�����'p�mbx��oB�����<z�$B���EB�&��l2cIn7	eJP�� ��8���5(���]���� ��f�y!�����e�l[b�Ae6��h�~��T�0�p2ϕܲ�n˰��	�kO	ã"sN0���"�ak���%�k����G(�ZV �f�q����`��>��܄��i|W�V���&�~C8@�
pXR��a�ݲ]{��8Y��)"�0$EL5P��$�&�"2�1ٵs�"�U���2�g�#"���jD�� 2���#4S��N	XQY]�G����9���D�!|GC���6$����:x��fe���8@vv�;	�݈�iC4��]C�#:�1��N+@dj�l�NHC@�~1v3�rXr&"R�n�1�H!�R!�Y��H�o����"(.��R�:-Ǻ��n���1&��O���
NP�]��3�f���$L��������0�N
K6�q�qi<6���{%'P��&�l�F���(¾5�u\d�� ��Bp� $0�����<��_�)��_��k$,+�a����FaI����e�`Z� �'C�O��\��~������Uݕ�a�B �ax��X��*�8/���3{�0�>��gʹŸ��߰m�b۸�ßI�(�������Q���q=ʍG	�ǎ��+����#>�у�4q _���?y��|_�'���w����&�aA���fz�X{e����#r��I ���$`��M mY�GA���<
�#{`����b�ۼ���v��.��~{v�F�}�|�<>�>��E�0����=l߱;�aJ��a���y��=�����O?���{�{��ص� ��`'�y�S���.l�~ �lߏW^�V���؏�A$sD_1	�_>��e�]�*�W�TJ�:I�R[V�ѺfD�>�EB��J>vG`ֽ|2�\��°@؈ l����a;�2���&��D���6Q��Q:�!��A^�r���!��O����",�a�J�O?]×#���%����O<�T\�X���g#�T^���h��'��,�� GJ 8ƻK,���7	�7� �ڙ�娞��3�2�)����*cK��um���*��6��!9V�"±�WV�0l���Q5�x,�y]��f�`���дq�����ќO�b��U���Q��z�����4��,c��l]l@�tp=r	��]�\ك���p���=������7���'�<�T(b�';�s�n�y��x��?�q:�~�����d�2�	I�10���O.CzV&
��PS[mr棷�۔a���DeE	@�P[���l�d:���,��ؓ:MAr���:,k��k��W��r�в���8>:���5���]�kd�]�xBo"��q�'�(����X��Ւ\4D�jKFxha�Y��hin�s�<���ß��g�3|�Yg�����_��/��٠�ۻO=�^z�e<�����{q�}Ķ�c��G�<�T��Gje?�8�J�%�����y�f��m�w����>|��#����g���׆�����\�����|�9��	v���U��
�7����h2V`�*��&��2U�R�. +臭iҺ��w�EL�`� Lk\���UzO	�u�O `i��#B�i���y,����r���]B&�#�� ��,������ы���pp��j�bSp���:�KT9&ٛ�~���n���n��8}T��ׅQᜏ�4��ΨC�K��l��s�¤p���(|�N��1��.E|n9U��B+��ԒH#��T�BB�L�U�Dl5����Ͽz:j��_tRj�;��L&�����	�Q�H$�ڲ��FTj�3�S���$:���|jVBc��&؍��&�xx|*bmH�-CVa5�]HI/BqU:�`�E��s���U��a�eX���Y��}ӑ�W��8F&!�oX���(DS��.^��ga�ʳ�t��c�/0�շs��]�DG�\y����U�8{liE�u"0"I�BD���g��?̆�tnK�>��v!.�����#L{���ÜQ��Bn2���+2���Ad�-��~�\M�V�L�g�>|oæ0!U��eQ&�8�aO.�_�U?�2�T�E<�����%����U�a���	�*���y����0�� ��E�"�����tT�Kg �}{,�К�Ÿ���G`������]��OV�{����}���{=t#0�����ǎ��$KG	�Gq��!�Ɏ�D_~��>y��*v�.aT�\+�ı/>ű��+��|s�?*�O	���6�y Y����qd�'H�J���,�_��`�1���-+XNY!���X���|wl�����cx��������a��"�|�nl'0�9����?��>�{���g���v.��� v8�w?�M��;��;��G;����G_�����㑧���KnBq�6D��!t΅�~�5l�j!����R�	�Mn5�0Ӕf°[�ʜ���#���a���
V�N�9��ݿ�_�In���p����(���10��i%���e�=<��\�\6��:h\%�Ux�8'V�yY���`�ҩ�܈�y�U7�\����|�6X KX�t��ax���d���2�[4e-�杇��k[1A��@�+�A~���P�:��,��}� ?� *��^!�X��jDu���*a��'aXeq7e�h_|��5o�a��h���M�`%�WV
�En$�m'����#����r3ﻉ ցrvfm�g�h�L������28��:�LA{G��084�\{��^,Y���S(��5���<��ÛW����r�e"//��5(.�7@\E��*E]u�������t�7� �%X�a�+E.V�a��Z,@�@�
rh^`l�Ĝ�F����p=�Q[Yl��L�]����d�R�$D��<˚l��^ӥ<�)��`É		�Ô�ɸ�����[�l1Au����U���	˖-3��/_�󶜇��n8ӲPX^���z�7���i2��\�mu3ȁ�����+7	�q�d�͋p�V�2(�X(;V������#�5s�������	�`��i�'T�.D
�=���MJ��1��s,vu�ER����ִ�?��Wb%���Pd�J�F�8B�6A�Ԃc����Q5���aDSqu��@�O�$°Wz/�Һ����mJb��7,׉��	>����Ϭ�0�A�F�8��+yJ/�Ôr��Ki����'tf��w*�����K1y���9�0��KVc��X��\,�|V�s!V�{!��s9�9�u�͆�b�s�T�x�y�;����o����Y��f�����yHo���ڹpTp��j���B���n�F����lGpL��(��#і���e���EKQPR����E�"#;)���|/�� gd!+��_c'�Θ�cVb��U^��Vm������.5R`mem�9HNM�2a�gr�[�������Ƴ/���b͆sx����`	�L���Ҫ�c㓝�����$�p0mKGD�	Ʉ{�}5���m�⽕���Ee�9y�i��*�ERFb	��|x���
��_[��v��!�i.��֣��v4�X�D���x��8�|�4��T8"Y����9�q�85/E�נ�y��^�3<��Re9��	�K�&�L����(��Os��L�1�C��.ƅ[���o������g,��>݃�;wsy�_�ae�8%k�Y)q���3SY�EЇ���'�b�g���ص�=�?|}�T�SƉc���������Wwv�:<
ò=�_�F!X>���c��%�0������0���F$�߰����S�{>y/<u7��N��̽x������������-P\WkF���
�TqZ�,�8i��p��Q���i+
�QN�-��EnY'J�9?������(n�WI�ŭ�n x�B^��B����Ѱ���[VR�^��x�ȼ�e5eʍ�	��	X%�����yN�N��/�& &�y�*��d'+����e7�l�}k��Afc���Fm���
vm����{�,"y���	�S�P�A����U� {%�~��>�T)�k]b)�W�#��� ��eNi��j��c%>Ӧ �
�*�!k�
\�7WE.��uS���%��Γ*�jc�h�p^�rv�����<F����*!N#+ϰ�"�WXsg&V`�:]K�%&���}��e�J�v��,J�?�Q���6�݄ W)~��|�0�'��	u���ODHX����Ͽ�~s��8c�xq9:>޾�&�.>)����F���c\%�l����4��*��	µ�zf3��E����全�(ByqaW>��ϰ��,@��V�Z'`�J��4����",˰�Y���!;C�v9��\��n@���mը�,AI^��;Rde�,�va�n���n30�������������"Q���N?�t��6!!!F���T7n�x��?�~w�x����A,�؉��":���3{��#U^�5n

��3ˁ`N7���iq�|F�k>@�]�n�JmFf�R�?g&�a���ޓk�K�|�5W1�|6c��d�/AV'���(�ENr*p���p��f[&��P���O� �#����03[�ģ0��b*�z�q	"���+c �>����4@S1���z.�۸�LJm�7!؇�K���?!X�a��5e�M!�
�X��K�5yϾ��G�������u�O��/��ԗ������8��Ǘ��P�~ ���5dT̅O|=ۨ��� %��҈��'(�pP�6I��D��c������ϡ��l���������>��{�|W^�s�584������Em�rw�c����z�j8.SJ<͕�S��N�$���;����p�"���`�s``(� ?���>�~���6qI�6�:�p��a�ylHN�@؞[R*�x��/ ��u[
�N���9o�-��c	�و�K��02����օɓ����	��3w��!�y��x����G���/��ǟ�[���>܉�� �py�EW�c�02���*���y�s_�R��l?g ��Ct~Xn��`��F!�b哖k��/B�|�	���a>���8��P�����U.B�2�jͯ�a��#�$N�� L��Y��D(��C�0|�w�>�g{?�`x����`d`�`�a�l`�}�C_���۱��w����/A��|{�3|sl��ۗ ,-�1
��˃���qy���n	�S�%�d��r;�z�z�v��p���ֲ��-�&����C���C���Ώ^���އ�	����#��?ނ�/��<�{�����i��I��ȑ�����"��;T���|�g�#�f�#�^��ۑ]3�tePх�V$� �e���Q�3�N���ִ -K��,'����eRS\�H�R	�r��,��1��ǖ;Q���A:^)��k���M��������u�0���f�n��m5;���f'��Op�3.
x+�XjM,�`�D�!&.�^G�c�)`�N)x.�b:R*�#�i!����p4�T����B�*W����
�s��I�VA0vqA�r��j �Nx��^���ka'x
b#�i�����2* %+�o,_� NkY�B�o0��%9��d��a8�0�ӵ�����eM�ۄ���4AsZ�޺����B`�R7�9�4j�+�N��g&U�ڸm�p<*u��f��0	U�d��{�c�ی��^�6t!-��U>����܊֎N�),/��,dp�Q�Ԅ���ef )������ k�l���d�$�KHW\��R�*�r�I	1�Hc�I(.��BUYʊUlC�sV�8Y�(�TWm�D��xY�H�u^�[�����U)gMu�RBp]U)�J���B����퍵T��5�"B��\�h'�[rp>�0��� �q��
�,�+�^z)�,Yb��W�3�exݺuX�`���F?������M ]tZ)RJ�P�>�����H����Hk]��"�ϛ��l1����rpW6��'���%��ä�F>�s��L�3�� <����H��e����+�|�z��g5�B�Qf�C�?>o^.v�
�����پi=���4�i�	��`x��0��jn-�]u�N�;Q�.�� �f��jY��6�30)s ^�aW�L%�� ��Ɩe�;g�o�1嬽�����;9 �$�X0l��{�jnlS�U!�SO�8��g�`������=��h;^}�-����&^{�������ӝ�t�g�����(�|�-��8�-�1s���Ŷ�׸��gu��>�]GH��,")����'����pBZ�ǥ��p%^���9����ؾg7�}�Y|��8r�|��{���q͕�ǃ�ރ�y�<�$�Oe����8����m���0��6nr�wBsfF��j99)YYY�-(5Վ��8��8�L'P�� ����T$lm	�׻�仛A@N幓M)���D�G�<7!�m���	
���/j�n�߸	��,g�PB(�A~~��:1g�|�|ӭ���?��W\��ބ�_y���{x��g��;��{�q�}�a�
�3|�br�a���$[���,�Kd	�Q���%�L�~]����2��-�r���O�J�f��%�#������΁�TS�F�a5O��3��v"�c�'Xn��^L^n`اr5A�0\N&{���V�c�`�������k���=�@�p��h�p��E8��kq���7�w�����vo߅��P��=��O��Z! �F�6q��9@0��u���������O?�'�������v�o���]8J���@�Ց��T|�E�#�d�4
�0h��=�!A�������=�>�y���x�dI�e���&�N.;?|р�ߎg����w�>�S/?��Y�pZX��J\���n�w#����B�;G@��m/��MN�|d7/0���2���EHo[Bx��eH�X��h92�V �m9!��C�Jj���!����1�V�
�=~£��ү�a{�[α�/L�37�
Z%��X^/��u�"Y�n�u��?�wo20�)��Q8͌�eݕ�V�me��QH(Tb�`�X~M)aY��
��0.�#�W�@"�k_u>�:B��عG�y�5��0!8��0\�)W�"r �_. V�4����І�3����detp��Cr�L�<4XJ$h�Ѕ*��<��A`U6A��*B8�
�;� ���%��`�(W
>�����,7V`Y�c�� ��E&ݚ��U&ZY#T��#!WE=<r4���$K��a�(':��~:?�f��\��{���6n��!�y�x�����ƭ�߁[���r+6���x^�|��'x���h�D'���X.���墠��f�L�p� %�㛫7ŤUS ]B\2����q&���&tURYY$$��`�F(�Zog���D(7q��&!��Y �Q��n,��5娭(Fa8�א�DUI>jˋ��m-u�h0���p"��9�0B�TtC������/�>��̜9����ǟ�3R���O`�6�_�<Oxy����}�=,�p!����`�]��g������
tu	�Cl�8����ZE9��n�8������So]�-�g2l�sx�w���|>����Y��3��:��7;�LP�y[5;�6�]�(:)l��SoD#��H >�GX�� ^=F�bkY�Gu�c��,#/CT�2DK5K�����֍ߥ��w�ƱU|�[�s @()�{+a�����0��P"+1�����T&Y$�b����ĸ*p�p������b�Ƴ��݇���F+V�Ƶ�^��l������K�������op�üu��7A��Jb��v`�Ln0�lM�B��]�s�hA��P*���jF6I�~�m����O��:>ص�=t?.��|\s��s��x�{p�U�՗_��_|	_  ��.f�c�O�XSmH�I@nFߗl�DF�F�b�F�-%q��pJ)+L
���a義�籲K��������o<�c	�R|����3P�܄s�;���&WVd�mT	���
&���Ӈ�cݚ���q�y�����a+�x�1�:�Tu��.iFhF�/�����MH�f�2�� IAY��e)+�5/�~l�X�G2M�}	�>|w�39��ub�G`8�������bS_�=�?�PD���\K�\C��0A����������Ҷ���5�U0<RtCZ�{涅��W8g�]*�`8�je���+�00|��7��jr������x'����t�ܱVaê���`���Gd����/p`�gطw'v���v|@ރ��G�܅#��8�_y�^Gi*��0lY�ÂY���Oև���v����#��+�\&��ˢlY����1��e���x�>w?�|�V<��-F�?�Q⃷��,�]X$��Ṗ�#h?E覷a|d)�ظ�fw#�#��ҩ�&d�CHk%��w��a'X�g�
8;��pu�BZ�j�a���0�l�:��d`��j_C�d&��0l26�=`*	T=2�J�Q�Z��y���#P��c� �x.�pj;!��É̕嶟#�A��"/!7#�Ph��T��d���2�0ATu��K<�m�����0<�",�)&H
�K-�-'�X0\! �b@X����H�jg!��i,��sM�gg�|d��m�Lc	��t˰R�	�yYs	��/b�hY��7(`��W�;�:!�%:�0,7�(nS%��`C9A�-�	�=r5��O�f� �M<n#ʺg�������>��o�7޸��� ߳�p���?�w=� �b�uG��w���cG��;oa�r s����t ő
�=� p}c*�*Q][�&vx�e�_����9(#t�����Gf�*��'8ŸJ�d�R�i�B'ð|�ۚ����c���X��S�	�i|����,^G��K�e�K��W[�y��4e���3�9����@��#--�t�w�y�i�w�؁�_~�{.@W�A�2K<��Cf��{�Gq������p���������K�Vކ��:�g8���(>q3���6
͝L �"@M�w��Z��]�T�gޱ0\6IU
Кn~�Pv�qv��zr�V!�Ӡ�.��г'����$Nϴ�"��[���ț�	�-VA��������Ws�Uc wT��q��.��Y�G���Q�K���o��tu��[�G�� �mt2�$0g�X��Hn�I��Q��8����Z�����u8��-���]&�����i�:u�ji3��#��4Q�� �[8�K�:~ן�_�0{�z�s@���9�Q)v�.�a��@��y�fptG8�5�鼚.4�MC��9�>*��EЌ1��ʢ��,.��,�?�9CӐ�p">���4��m��&#'-�q����4�9]�z�, >AZgI <V��!xT��0�s[0́3�t �g����Lt������Q�f`�}�x���DCC1upӦahp*�
�a�g��=���*��J@��W��� ������Q��G!9
4������XүJ������_�Jm4`l����e���X6���/ۂa/7G�/䳼a�R%�&�b�*��Lu�_��D�pD�2W�D aػ|5&���������X��/�����n����� s0)�� g�U�N0��ۄ�=�a�G�������oJ�y���R0|�0, ���C��a��ػg;��r���w�T�c{�珩�r�C(�tj�,ˮ,�#:�1��G�1ϯu��ˏX@|D(�tlҟ�V��]����x��mx�����=[�����Ͼ��G�+���)00�ю	1e%ǜ����vi�Z�Ԏ%�2j9��Ni%����.��I�ax�\\g�M�$��@��A�$<��"�ѯ�a��Uj3A�t2��0��<0l�X�!ЧP6�=�.O�\K�k�����60��wRة��	��i�H�DŔ�(�^B�m6y��ʦY����$����g#���L�b&n_�Q0L�(�eX0�)A��q�V�n�@,% �aY�)��
�c�e�r:�*f�հ i���*���NP,w	e��q�Gy�x����Dbͩa8�m���r �UН�����F�b�l
z��X@le��x��x����*��~5��i�#��_v��#n�=w �U���*�����^gz��s�,� ,:م��&���l(��s�*�޸�]�Hv�as�"9����c 8-C��<�VM�&�
	��H'rs�QWW����:k���i3��U}N�1��At�^�W�K�Ù�e�U6	��o��V
5�5��.����j�b�y��#�iY�ťEy&��@�fK ܳ����á�������<<<���^�^^^����ǿ5����lTUU#�f���l�N�@lZ!��P�寍�i�{aU��,�J�v��BV�J����) ���e��>v�a|��%bRj=�L�2����@ҵ�E��ϣ2�p:���}����yJU���p��w�0����Q0^g��@W��0L��g<�[, *��AĲ{e�!(��l�	ı�sM�	���KQ�������o	�Ä_�W俶y�	��`ɲU�N~��g��҆��g�=g�\}�58��r� f@���[�Gc}��ͽl�*��� �vsWmD|^z���տ�<���Yl;L^u?°��A�'�p$AL0,W?��4������Hxx��gbcB�_|�2��-6�'a�ig"��[� �c��hGb!6>����`�`$�&�#�AH�������$
�l�H��Ʉ�$x�k�Q��ݐ�0�9iۘH$�m���ߞq:|�Ox.-/CFf&

���n/���������p���"2%�uU �U��,~oy��Puڌ[�~��,qd��k���	����l�9{I�a°7��`�~���&�t�kõl�N������UOt��`�����^�a�J�p�L�Y0��� �pD�J���37��h>۵�0����j>,����	����g��o�N<�ǎ������W��+N�!"�GP�H��w��[U��&g�;P������]�?*��1��\'���s䐶�0.�-�K��u���>"s��÷�6 ��]��A��{+�x�.<����>h`8(�
~�| ��P4 �ۜ[>jf��Z>9�Ä��Ji�ZD�\B-���NN%;V-�e�%�K�a�r�8���.�ץ��n���Q'Ept��WaX�y{d,�#�]�[#�kx�5�Q�����D��I�>��J��!���S��)�,�	öz�j�T��V��nj�4T��0I�'*��ӱ0쬙cR�	��z�d�k[��
�iET~��BN�-Ŗ�׋ز>#�,ı���r�*D<_f�q��veS�XFȕ�a8\��q��FEB�	4	�_�I�2l�p���;V� :��Vc1��`X�aog��vn7h��G�&�*���枂�dA���J�����`>�� T�C$�3�%�_�@k�9�V5�Ͻ���l3����8ܰ!,<�1q
�h&��c��N�8��"�.�A���ON2��vG���
t�$QNp���`�����p6;lY��J	�%�W��C�qI^�V�@KC��\��\!d�-�TVb�O�uB�崏|�����W	��e��0ǸB��[�yA�\&�J���|����V�f��l����y��� ������ʩ����0�`�@��`X��T�#88��)�Ą	M5��H��E#"Ʌ��L�fU".�!�|�Z�I�#��-",w�ɀ����3;y]��(%�~��$[ۺD�)�H'�f�!pr@vFb���ܓ�gq@��Vn&���pZ#Ng=��[�o�s�;y=��m6���f�p���
�m�6��v��6@,˰�ؒ�����\�u�L�@Z���D@<g:�11����o�N���ꆑ��Nv���!,S�����wC��69�Pz;���i�ʵ��{�~<����68�/ƶ[o3%�/>�"|��{x�ױy�&>ו&Hm����s�v�?��/B|n�	��h�c�"Bs�N˰A-�
JmE��� ql��B1"e�v!ܖ� �mTR"�8`K�p��8�TQ�h�G]E���8�#"	��H'��fd�es !��t\2�N� :"��H��99����US=Ӫ��y�7멤�D�-�p�&q*�Sr��aB����#�1�k��	�^���e`X�8�vd�䠥���������jG.��m������{d���pTZ9���S��0SR�)e�����zc�կ)2��(�v�	B-�]k�(�Sd���ǺJ��t��-|�(�l�39�q��e؂ᰪ��f{|�`�N��%�٭^���Մ�u��5n^��`�@z2 & {�_���eOG�eX0|j��%y��F��$�6ػw7v�ށ/��|�%���(Ov�~s�|}�0��P��;��:�?}}��?}u��o��y
l(װ\�ʽAiَ��w�|n��5����KY�wS<��>���/��~|wl���lY���!����2,7���z�mx�'��㌨X���+�	zT2^�:L��@���̺y&8�IN즺��EH"�$<����V�V�	�n��䛫�4��^�D0��ج;Q.��_g'a�-W�&�0��������j�~��ֲ�(�u5�(�$H�Ŗd5&�3�@�R�iY2@�� �}r�΅�v	�s	��n
�M��t�_��Z�3�F&*O�ՔX� lca�v�Z-��`ʑ}Jŉ0�ۺ�l��{,��&�Ft"���Ԉ������c$��A�X��l8��<� M8.�5�!�y�������z���C���8³|��a���<>Gȅ�p5�ag�f,�r�p�,`�c�E���B�"�#�A^X~�)�����
��Y�紏�)j:�j�Qr�,j�	��4�\�N�T9�� ¨�fd����*L���gchh6&O����?eC�g�o�T�N����,X��,�����ւ�;%�be�W�T���ѝU"e����2ةU!+3���*�DEyʊ�Lj5�H�!�
de�U���EB�`A�`X�H'ؕ̲��cI�h{b,�x|cujJ���g��������rB�2N�e!�l�'"���p��ADpH�����Æp�u����֭[�X �tZ?�^r�%���q���c� �h?��˰t�F,Y�f���"u��VJY�!$����n��p 6y�|/kkqp&�I'���/�#�;Nӳ��/������~��a�Hx��d1��m9Њ�����Մa�;m�[�q�K	�T��9^�H�����%Y���VbԎ�្g��5lW��#>�bBZ?&��)�������|���`���1�p,%ZMKFdoXd�޶�,�U�a���a����Oc���L�y看eKW���������3�#5ŎI�|�.�����c�o���Kb�Ct��87�8�-��6b������w��4��bE�q�ДJ��``�j,^���9g_x!6lވiӧ����-�koE'��|�:��сֆFHR&*>*�1��hBit�bb�b)��s�)���PUE��W�We�(��O"<�X����'+��%[ �d�Y�,6P���8*� ���(�pp\_�<�8��=Dp}n^�ϟoU5]�AȕW��\}-���ո��;0w�ձ�ȭC�\$���>4ϸ7??o<L��4�At˰]~��j��a�~֯-��d�p
�=0�l���U�Ye�-��7�>a�����ȺE��xx�<�d�`5��|��E���G^A^I^C^O�\K^����p�"j���P4��-����&�gX0|�{|��c}�Ga�(�� 8p����;>�'�|ċ����Ñ/��;y��y�/q���������:�G����;�8򹬸�@�U�N��ZY)����˃;�{���໯�  �|F���=���M�c`���nq�߿?���sD������kn����x�����[/b֊%�JJA`n���[�@e+9L�F$�x�I\n/2�#�s��{�EH�^L0^�$�p7a�k�s�X��Z�6``XSY�	�i�����Y瑖=0���_� ��pj��-{�F�kD0�Ir��y-�	�Rʏ`x�\�;>5��(�_�7�Br�*$Q�����V������'�IF����J�e��R�\/r�6#�v��z��QR2��Io������t�&��X�	����YMQ��mus�c�U�l�O���E��6��"����% �)"S1�w�*�[N0�b�TnSF`�c�c�ÄQxN�b�-��M! �B�5d�h�*�N�-��� ˎ.���2�"°�q6��[M�5��R�ŔM!����*;��iR������g?mW6	ApJ!ǝXh�d��2D�K�O�Y�)�u�Q&3
��[9��7��Z���~o}��=�nf��Ï�7��ͷm�}=�}[.��>�G��|?>;����}l:w�q�H��KN�`�0��E�%H��4���&$�"��\T�O�$h�$���)U�FK�L��L'�����������|�V��$c%V
��L�q���X.
����0��:�@��Pc2H?aq5�)�pmE����T�}�"���c]ic�6Rt���y������o�>4'���7$�{�=�ڵ/��z�a���>��^~w>�4�݂��f9����w��#g����3�B%��10l�]���n��P�m��3���v����pj=;v��m��nۛE���l)%T0���F>?=����v�u)ؑGU�?��c���0e�0��@lA�s�B�M�$��,��D�W?�e��"��\I �ߘDJ"�J	����$U�Eze?ν�J����)��j�2��i=��V<��cx��W���/��������{a��,�9p�0�o���HN,j��n���FЎ�=ŖNg��l�$S�R���3`W�~�)l�n���>���>ڻؿ�ػ=|?��v����x���p��7bӚU��������o@gk�Q1��87�����~�����6JN6V�D��$���]3 l�y`XV�S��o` &�x����y�}�SPZYWF:C���{{�@�
B�b��X>��Sx����o������[�����E���H*RJ��^(�~�3m7��bNKW1�X��
1>ٲOL����W�Be�u���0��0�Ɂ������W�	��R�0�^?��&�	���FV�D�����@���)�����շ�o�����0,���'�,>f����#8��!|��~�޽۷Bm7�l�^��ڋx��?����qU�����W8�o'^{�I<x����K�K��q#��+p�k����'��ۯ=���cC��=x��mx���k�{����x�1��o�	w�q3�����x����7�oƓ�(S�]|y-����J�����.X�K�[�Kݺ��ո��K���bå 8-Q�Plm�߶ �|4����qd�f`8!�Y���%��a��J�߻��K�Ի�=+`�^I�"x�b��=�{U0�E�MsK�b�_�5/���u_�p�F�=��30���ݚb����p�ey�5�yM��°���y̿C@��)@X{,�# L%Q��a�Òa^'�m=�W�`�	Igi�#m��Z��~�S`An?T*5������S׏X��f�s�|f٠e5��ri��L�_�r��u
ބbʀp	���nB���#�MX�t�"S&w0AT`.�sW�XGdw���}
��U;��"�P2��~��&��b°�a6A�T�,���kf�:�&ݚ�W�6�'��%X�a�_���&<P�˟9Q.#F��,k��"<��g!�b��7���߂���Xv6.��6,Y���-�9眏��Ƽ��8��p����ڍ���SO��7��]�߇����lIHLa��r���$Lэ�bK�ܼdf��� \RR�T�f�3��I�$��M!?��a\%�)�-����R��7u^����T�Y��f�	�kςc'�Ӗ�b+7	Y�s3�ʍ璋D�ҩe /˅�l��WV`�	��=:])�X�l����i�����ؽ뮻0u�ԑ���Ӯ���x㍸��+q�[q�Y�`��L���s��}2bs��*CxN#�s�+�'����O)����l������!�C�>4�� �k\'R�����g�Ϣ;�@v�!��g�ޱ�y�&�' [������`��կx>�M��а��F|��$�*���������a	��0!m �]����p�0ٸF(8N`�������X�:Y��U���}^�n�|�/��n�n+�{�a������N�� >~�}\t�9hoi@fF||��;��>؍�_��Vm��Ɉ̪�����vC�I��7`\]�x_�TL>�*���	a�Fn\���w?�y�E����x�'�^��n����������b����?���}��W^�̩l���JCBA�$���1 ,k��_��=B%ǫ��P[[k����9p�7)��c�ux�<��a� ,�����_P �����9����8	�T+����z�����3�{�?��c���{q���'�õ7ߍ^����^���������l'��C�,U�Q �>Cm�\�|�m�'ٛ�}��7�l���;�+�ԤV��Q3���30܋�)��0�w5�\�Ֆ#�j�*����-T6	���o��w��xw,���&�u� ,_�C�޳w/v����<t;��ă=�k��
�?�/B��w���� a��'�uW]�e�`�� {�0��C��;�ˆgb��a\�e=�ް��-Ċ%�q�e�W^�c=��Ӧ"?'�E�b�X_��*�4[�j�C_W#�:)N{;��Z���|d:��JB~��vv�)��K����x��l8���4ySW!kp�z����d�#�0�T8��慦�Aj�"�*ܳ�=K��#�$|��	�R��rj�ZOE7Y��i�b#Y��
!YdcE��aY{�c���y����vK��M��ݭ�o��y�d�˒�~`Y��^��ߛҺ��U�A�&�U$E�ANV����Qr�r$5����1&6/CR�rB�
c%N$<'���6��`��l��v�,�D~>�=��zV#��qt��ӗ[@\�v�ӑ׹�CP �l%t �DV�(����VеUS7"���F������|ْ���P9e�;�8+߰�/˺, �*�D,;���.vHTY'��S*�����bn/��r?MU�c�T6`Y��i��j��.��/�pK�O.���b��FBi?2[梈.Ax��ο5�g)R�f�?��)a8���|�S��n�%S�����"�&��8����L`���dI4At�(Y�w�x��u�� �t��f��ZV����/.�qN�F!88v�Q1��FLB"��C0��!�(*+G{w7�	���Uؕ��T�$��	��r�a�KT�� ���2a�� ϤXS��R�kC}�q�()�!����YyK�
��Q"62ԸJ�6�?aA�'��*�)�N��e�mA�\(dE�zmd7T�W�R�g�s�\S�#��e�\��Oe�]�qХ�&��PV	��
��\ÿ�Ϳ�Q]]��:�SZ���y~Nּ�B?3��*Z�����X���\��ʪ �V#"We�;�ϰ���aT�7�l��&V}]ʉ��2���C���{OQ*=yo�A�^��+C�����G0k�E�U�`���������K߸���g`���@���>��'��/Q�d ��fG5r�Sh�~'˪n�aOʵ��.�E�Ĵ&ß��wZ'&:Z1�ބq�q�uƗT��&�6c�� ��@5���l�C��X��|l��9^}�l��F���c��������Ce=z�n\�ɽ|~r1�����p���؟�7g�פDd�"�a߽~c�(���7�Tn�*���������s�bRTb�J�_݂��Θ���.�r����4�r;߇ƚJ��[�x��kV,��@?�	|�b����.��jTd�1bCs�j�p!����T[���CKS3�%���);%K��� [R�
ɀ0'������ٙ�24ոT��>x�!�H砢���f�BOO���իV�ҋ/����r�:\���t�fT� 2�>I�M���_�ﮖ�3>�Vna�=(pߵ~��0�|�eArl��V��}'�LW�l�Ҫ�Q<6��u���ܖa�,�!�C�2Q��U^1�|��������\�Y� �UX�$|��`�	>�+�b��ބPÜ���yd��^���ħ։���~%q�0���s�<�/�N�� ~�!쟣	���8��?`��a�-��7�2�$>�p���Ma���~�Ź������d�Q�a�Ib?>#q��s���3<|_P�?��x�W���_��|��q|��q|y� ��>�s.�pAwΝ���'c��iX�p6�/��K`���X�j.�����Q�/?�<�~�V�b��X�p!V�^�u�S�v�j�Y�
kV��V`-��֯��u�v�J��"�Y��߈-6a��5���Ǳ��9o���Z� �9�{�#�j:��ЀX>�I&[�d�#����/FR���2�k�e	6�^c�ڽ������ݓ�� [�_��a��lD��h�)��@�fB�f^o�z6�7���&�n�4%����E"� ��&�%���P;Fv�k
!V���ɍKakU���}�&7�sl����1�q�[�sp�EP�I�k	��MHh%���7~7#��밤�D�s�����'h7�E �1 ��%����#��؄����>l��)g�23ȍ"���׹���E���Qؽ�X�4葅%�b*2��|p�)���yڐ߰|x��"� ���nbI7��
�BE'R*9��8p"�g7 ����=\�O��![J.�C;���yH���8�udNb	�Q��q�D�Mpv"�q&r�o"�:���5CHk�{�R�uk�|�4�L�UU�T�~�."��@�g"�v6�j�`�A��8vn���9�5�Z�	�Ӽ �m�c�e<����ΒF�r+�Hχ+-��ZB�̓�i�=���r�`�Õ���B��FF�)����a�0;2����
W���������4d&�����p;s�)�D�3���v�5!��,ح�P��X������^�A�Ȇ�W>�r��*+6˞@:А������v�Jv���X��몌���F�h��ْT�9�~��3NCLl4ZZ�M5�_�E��UFE�5���
�Sխ��,82��VXGA9�K�Q���y�΢��z`X �-� m��V��DNk7���Y��B�|Vl��� ��f���w�Ͻ�z2���m��#w��͘�i��.��m)��aB0Ӱ�G7.Gd�rDP����?����:�k�@��#�)��S�U؇ 2QV���M�L�aS���$��g�#(�ضh�,zA��X��"���^x�U���l������-��;\����	��~>֮����F�fec�D?�#�x��A&/�?zE!��ｸ�W	�=��5U WT��A���'�W��V���f�؋��wx��#*�^T��싘� >�Xef��6���%^�0�c8(�6!6�Xu㤸8�.���P>�)����pd�9���@5k� ���M����2e�K�7<R���{�,�c%���Ct\,�u*��ɉ�^��z��4���;�4�?��-k��|��ʒ��i,��l��"0 �����
��8�G;�A}ln#�y«K ,5P�~��L���0��0����Z,W#���n��`*�I�g��\!���%í|������'������	�#��ӊ��{<�ߧ��79���xL����W�^N^M��@X�$&�+ϰ`�ĄQAo咟��9X�s�k$^L^��������i�_`*f ��UL�4TN]�-W_��Ӕc~��7�w�>|��'�����j�a�*�S0,�s=�a�Pt��"�ai,�� S������,���}�n݊�^{���y�:����O�ӟ���W<�|�������m�Õ��͛����=�l\x�����x����/c�g���٧�ǂ��q�Y��ɧ_��o��7��o���ڍ7�ۉ��َ�����>�>�{�»���饷�2����}���+���W?����C�����kgA� �&7#�r;�v���9q�&�r�ý+��+h� HN1a�5�DN�^�T7;�3@��l�m�`XPl X������,�b�U�۲
�U*���%�-�߭0�tg��6�����ep4/A*!��4�q�R�{:Fvv�'���8�f��s��N 6�ܲ
��`�H��dq���@��2l�'��G�ԍ��[�x�Y-�C�.��y.�	���7"�c�v��6H����h�w�Q�-(����РG	)53HWO#t��������v� ��D�����=��)e-#���b��*GTv-
�����4rچ��^$�#���U?-3M��\l��5�N���r��\܉���o��$Bt4a8��IUS�h��4B�2DxJ7��oJ����9~U6W�sUL �g;�jlus�=͇}���|3�K�斧��G��-$ls��9���2��މ[�}Wm�^t.��RS<`嚵����qյ[�t�J�:q�����G�w݅��M��i��&���q��9�2	��1\[]���t��c�Ω\z:Z���i|c#�5����X�ۛ��'c���*Сu:F��O�W3\��J��a��N���B�PU�֦z�0���
�3��*4F�����7��c�e�9����Lc��+�(�O�J�`�g�}o���14\��+q��7�[n��>��{��FdV9��[;WG���%��p`���>g��paX%��-�tÊ�K
�	d�mS!��aӁ�U�F�춪����RJ5BBPn�I����\$±lbe���p�`xa�@L�õ��=]�*uQ��w�&�w��V�fk���3R1�P�E��f� Mb;a��	|2���.xn���S�O>���ظzV͛���N�M�f��K�-��`V'jJ	���s�p׃����>D��L�NC���i�0���� �ٱ��%���C��0n��G�W�q�9�Ȯw�ӤV��9	�	�%[~�)�1 &w��"��mI�f�����o<��5��,˰������+����Ӌ:������srM^���h�#0LV�5��d60́b,��`�?0	�1���(x�x��3τ���y���Y�r@�����y�ؘ8D��sDB����8��	[1\z�� R�����c���@(a�n7��)��`98�Q%�쟦�\���>S��?���������c������ß�Iv7�-����%�Xb`���1��BV��7�}'n�}^y���mY�w}��F,�'kũ`X�����ϱc�N��lv�ۃ��� ���j���8��Wسo���O8��78z�k|���p�[9z�w�"������_x	O=��|�Y<���x��	ٟ������ۿ����x�y������	���a�E�ǅW܆�/��]~7ν�Nl�dξ�Vl��n�g]p=6l��6^�%��â��`����v�Ŝ?�6^���/��b2\����E�m"�6/Eb�|v$�����}p���m_�ܾ�M�G���	��a{��'j-5��7)/p:��hVZ4B���H�[��@��`�;��H��l� �0ie� ���� �ں��J�u��U�����4l�-���T�W�<���D`r5-d��
�b'��g
�R�'��AHv4s`��{i^O@�H8��8�MP�v��4ok[��pz�B�v# ���P��,p%!�E8��I)��ɦı/G�y�(�[������{q�sIC�Ѕ�I�����P��$�g���L��,6��%ȏ7��9��
�d� *���Z����9����t$� �Y���J؊	�E�f�U���p��#���y��Ψ4���Z�fV!.�C����S?���YH.��r��.�+,�b;�[����+�
%DOF�|�\�@��mTVWc����|��.��z��W�����ټn?�ը蟏��=�G_xw=�8n��v�x㭸��q�%����_4��]l��Cl�ض���;^���#��
'+�AXVaA�X.�,GiY�Q�<�Օ��h+��Vn����BsC�;�Z��؋�Z-�d��V��Xe�����_Ω2�����)�JV�m�a�|���F]�)Y��������0���z�	���?|o
o�_���e��^�z�a�f��y�9<��Ӹ��{p��O��ǟż��!����Z�A�숳�*я����ɈV����N�ږ���G�gu#�ψ��gj�Bә��J�o���R�A9�>������0�����="��j�UX9�	�a��w��H7G��%QⰊ�P�K~�^Y}���ӛ�Ӌ ������fw���_~��>N�j:0m�L�9�sf�Ջ��5s���x���n
fMmBQn�#"����X:�b�0�����p �e�&D��*��߷I�J�8*�]0h�� ~�^I����v�95]螾 k6��MgoƊeK0��mM��no��D6s`��K���9�,/�󜌰�PD`��%��c	�qTB\AX�"��;�|O��bd�g˯Ӯ���|9����F�*<~�1�%�	)�����B�1n��C�_�䇯{T*Bݗ�Q�nef�����CX�p�6l���l������[.��+P�؇��&c��d/�aU�"���T�I��g]V`�C�ۄ�JG�T=��s�%�th��a�!��I5|w�~�����~��q�(���J�we��0Ay�F�
ҋ.���b�/�����m��g��������y�}��w��ν{���:��!\u�ux�����'�൷��燎`�C��������$(8�w���������d���h�>�����G;���Z ��~����N�@�#���_;�B6���9��k�����ȫ�����ȭ����YH/�El�"��yMH+l���FI���CZ�L�!��!�e�Mm^Ɨ�a|X٘��I8+�!�c1r��J0,�p�r��
jRz֎ѺQ���f�j$�0���'�����,���
��#l�d0v���-��	�kW1g�*J�<�kYl��
\U^�ArzӚ�"�5�A��*��2r�R͌�VO7�S)|`�{��w�I3x<��!�U�^��5ƚV���y��p��C:���m*��נh2���K#�+����|�"�e� � �X6��9�^������	S��tiJ�6hJ8�/8�G�|�cRb&���9+'�E� �ل��Ĳ�h������?g	f,]�Y�נw�B��Gu�X��i�>u�j�La{���:$�T �������/�����U�\��/ǲ�.�ܕ�`��M��r3�,X�ڞY�윃��!�G'"rZ�FZ	�C�1E����Α�`½��=ЛT3��:	��D�*����<�hY.�N�*�!��3�M8�z)��%���4��^���J����B]Kj�ZPS]���^�kf͙K����Z����s��y�_��s����ˎ�%�6��X��J�/_a%���~��Fy��pN��L��3,_]�>�f	~3G X�[E ��gWY~=���?,ɟX��%�(%,k?ڥ�:���Ze��k�*PUYF�Dᡶ��U�,� ��5��a8"<��Xʁ�| ��aW�5e��ϰ:���rL�6S�L��� fϙ���)(�gX�ϵ�g
۽.Ñ���i䴓�#+]��1y���y���6v�.�pZ�#~�
 #�)� �R{�B��{'��':����td�2L���BV�h�í��a�@8�qax�M"�0��)���F�x�	�����PQe3���A��]��"��"��#.s]D�lD��Ct�<DV�ြ����JL�=5��p��5�z�"\�j�����6a�P���а��I�BBZ	������lR8�	�����!n���S��_��
���!�7 2�S�m�-=��َ�>م����{�p�z�-���M��sO?��W]��sgᒋ��=wm�M7^�ޞN��D"2*��O��B�W�b��ʕ"�JP ]|!��k%z��QW]c�X.r�P`����`��>�\/4 ��㻚�k�������hʳ~�ˑ���3�؂������6V`Y�u_��-7���:�6mE�p���p߷'�x
/��*�|�e�tǃ�|�\�>���P�8��e�V �Mb*bJF]��sT�ة��l��ڗ��w�U�� 5X���,�,�.­[b�2�"T����%  ��IDAT��QM�FX�<dMf;�B5��@��e�p�e,�ex�r���I`�JIl���y0l���ao��> �/�N����WZR�I�g��w�a`Xn��%���|��?�={��uB�_XV��c�����O��+���\�kn�W^w��e���6\��&\r��r��8�kpΥWᬋ���K���զ���ĺ-�s�Uf�d�yX��<�ނ��V��e
���]�i���ɛ��Q�/��zD��נ�{5rۖ�b2�n6B�f+���>�*� ��\ӷ
�MW���=���ٵ�}[�h^����s�^��0<d`8g`%�v��+l3 l�H� �=���^�R{�"�J�h�����0r����s����sћ��ٌ4n� g�3x�w��ѽ�]J߶i-+�jYJ�%�6z	G���a����NeU��x�UR	G�TbQ��]M,�2 �߁��FDdHF��'*,�~DZ�7�1�͈�nDXz=�	��!6.A;��F~�u��=�CA��5�~1����H�[H8]�x6��v��Il�ll��|Q��]�ˢ�wZ�����3:̠���[�>��謜�G�iMHf�Wй%]�ચ[�T��B��j��c�u
�Ay�d\s�x�����;������x����{P��������źs.��Z��3��/�3���臞z������}���#���/��G���;���/���=�"��u%J��!���ф����?{�չ�����3����s�{ۘ(	�K���*�s�BH  !���`lp '�'08b���cr������+	d��{���{��}a�c�Z��JU�Ϝk~s"B���n����N��e���^�_sO���3l��:����s���`)�A��* ��ݠ�4�� �e1�,L)gK�M�����p���c�7�.~~���"�3�^^�0�M<�Q�/����g�˥b�%Y�,�1�M�K�����8���@�P�mtd����'6��k��Dj��;,��$]�T�ϰ�pAUR�Iܰ@��
A�d��
Y4' ,�ɾx�%n�ʭA�^��I OIJDfz*����HC�j5�c��$���������?��QVR�tN��(��R�N���"�q`�}�pC���$,��4�I��5��<�$F>�0, ,�p��� *�N°U`�X��m�����t��J�L�Txs���#��k	�m*fX�$<̅l4Ȥ_�x��`�/�Ah�H�#³�m0!ح����
��C A#�@�?S}���A�k'y`�
�%�J� ���3��8���:���k�cJ[�^2�{�N��y�naV..���@���GX�O�~1�2e �^�k'����,Y�K���/��m+H�L&�U��K���'�������n������������#xe�sص�9<t���?�;���O/]�GDOO7b4BTt8a8!��/�5$�½�M<���A	𦥤���	��ZBqyiL���Z�0�nMB0ě+�R�Q�P��H�
�&�#%=^>�
�G���տ���k׭äɓU�i1(Ǐ�^�j�*,_�sf�ƺ;�b��7��GŖ'��ÏoÝ<�	�+Tj�P�^�,��_��Agdl�1RJ7���0��7Q�b��q) �9����%�xH�ȣy���|߬n��	'w��ބq�2���z���p/�{1>�^��s	�s0*c �	��?�N3V��C�!�v<���iS0�Վ���ix��!��{Fc7�y'�l����y�'�����/&?�?��9��p[�	�.�s0�o -����}�[:PT߆��f$���W����Ӌ`K+�
aM-�%%�*@\F)����3��B$'Y���R��at!!����W�r$�-��e	�M��lX�䪟�b��yLn��� �l��̉��OA:'�t�jj�B�a�l!!l���gCʓ�ˠ!k9��3LX�k�u��R�ոa8vH��9�p,aح��"��:~�*/��hp��!�� ,_��\]�b��R��~>L��y�\��f�D��RB]IL� q��NyE�ضB���"��lb%�b�s�φ�>�� I@����e�_��A<~�t�S㣓�CiR%�n��$]'�1�D���~i|�C������I�N��fN�����>Ĉ�V�Jc/��:DH�K��k�$�!��S����	Y��'��Za�i��P-���uL��9����pu!��/������0�#����������ip�u�Y�K�������������#�c����ؙS�������兝����ob�뻱��70g�RX��#�qk�OD{�t���u���}�ȭx&;�s?á�N`߻q��'���?�<�
�[�(�$�0N�����ZU�9���&���Ɉ"�8��ܲ����ө$5����P�R��C�4Ua�!�*2(9O�K�0"C*�U(6fW�UT����׶���%%hhhFiY�Z�PVQ���,d�䡹��MM(��D�`^P[�Cy���v��,Y�j�xI�����,2�<AW�Kܰ�,��#/;RNB%2y\�X����a(X`ؽ8N�`�J�9*!�%��(7K-��xb����51�x(Qq��[�����$�	��ٙ*�Y����~��p==<PZR�6>�u2�O��&r�KJ���>,\�P��"HT�����%H)�����m�\�IK�� g��i�0��]MP�	L	�s`)���[�bJ�9�?��30��>HV�a����^� U ���a��Y�F�nQ`n/��ֵ����]���$(�θ��<��s\������@i�Bo3�Z:w��U���
���=��~!�nh�)���k0�(���t��f�fU�� I�^�o���T�ݠP�m���0eV�fR?Z�������U����b4֖�@�f$!O�,��͜�����~�u:�|i���X���"#ÕwX V��`\�K����,T��#'+[y��22Ṵ�H�Vo��.��2����Mb��v�2�Si0���#�`�������#T���3f���J�t����aY�* -�&���ݸe�
U�k��_���o�rT�M�5��3l�a_���4il��J(�PYz���#���g\�@Y����
5�z���3W��Df��a�� <(�K��h�N^3�p�����H���i�X��ث0,aWc�ǋg� ���&����	�^O��8��G:a8�0�Ь��r��pF�T���=:��]T0|��)\8�w�Ꮞ����ŹK���m�cb�tԷw�����ې[׊��&��5"���	ә_;pKz	̔)��*�-�	���f�ÐTsZ9�,T&��e��b��+��E˲����07��X7FB��z6!RJ ς�eb
{0�^��F6Ɖ���0�jO��O�	�.B��ll���^	C�N&�a6xM|5a��Ʉk0\#6(°J�6�5�n��c�kA[���-F?/�J
`rk��ҰB�\���e꘩���x��.	Ã�aB��l�9Her�͜�ЌnD�O��P]��:͆-��JK���(��,'LJy�"��*�Xsl�B���!���`m�RPl
4I �r�A"H�B�9���z�uI6� ���2�,D�3�D۲nJW���"���5���݈/�[�T$�*	�<�/9<%��Q �	���K��0G-��@�1�%c��ۋ]N�/���t��¸�xC����f�ˡ6�ះ��
�,#��=
��5Ч�+#�א�������	q3p����ٗ�o�F�͚��.��%���֌�Z�mm���GCS3�/z���8�.h�c�-+���;1g����ǭ�nW��;�X�Y�fc#�[�-����7��0�PR���R05�b��@����7��\�H��X<�|N����n�,%ӕ�X��u���c���wk
�?^���I��"p'� �e�my��ڋ��îWv㥗v��{p���g���;p�;p߃a���	����۱h)���D�*)&6V�J�pbR�*�����&��4��x_�\lJ��­�d���v�93�aѣ8?[�JHL���pw�v)o��,��XΓ4jJ!7$<B^'Y(d��A�Q@,�����c���k%�W�W4���*S��p�Wb.}�Q���j��ꖰ��7o8��q�����̳x��K/cۮ���k{�i��^���x[rT̰xm�C�G�KR6�/I|���l��9�Kx��p���a'������j���S�%{°_iO�C�����Kx��.s�O��o��ܟ�*}���a�����&�>��G�n����$m���s��@���c9��;)��`ך�I^�ta���k'O��m��RD�V��"aBPLܠg8A�p����L�C<,E����+����}x�<,��*�c����x��1�F!44�����`��P�i$�x�~�v���`��Ju�Jx�,���˲?,�W����x%,����%,�����"�4K8�a�%��P�4�<�AB§R8H�q�!c���<�{a����(��7ܠ�#���Y�.I�E�����Y���/o?Dh�48�ft�l��FŤ`�.�LE��.)դ��;��[�5�Z��B��lDL�:.w�"2��Z�d��+�x�e�pV���0�ݍP�����O%;���e��x�d�P0<�0L�9>Mb�%Lb�
��ч�l�c�
?����?�3�����;����`x��፛7c�;�*ϰ�I�Maxx��YЧΞ��K�p�+x�7�:e&r+Z�S)q��p5"����J�d9U��*�2*�K)��2��A�\B�cBpZ%�+�&���*_�(Z���*�8<�Q���
���ڼ ֦��J���ṪЅ�b6ax94_O�$E�A��X�����H�[����H�\@8X!�V�6B�N���zr �M��v�;qMs�°�IH��X~��D�7X[�:�_���~)��+x|��X�jpf�7���i,u��yjQ��Tr�J&�Hu:k�\ث���T�ϐ�	���"�)��Tl��I���N��ܺS���
��Ct�F���@�'��	���Pa�TD�RaJ,D�!	��,r��3ʘ�Xk*��th,)��c-�Q��,��[��1:kr�`�c["tV,	i0ť@c����B�ͅp�y>>��t82ʐZ� Wv5��k��Kc)��$Z�Nĸ$cC#|M4�2Z�E��Q0Q��*`D�T�uT�_O��+AQ� *:破���AA��
i�G��wd"��G1�i��w	"��Ǧ!.�	Mӗ��g%��i��H�`K,���uM]8y�2><z���gr<V�^�Uw���E�0sV���&�(�vG�R8��� � &�M��g�b��E������˱}�v�Y�F�n�Њ���?��M�^EF�4z�ny�Q���&:4x[��8B<�@+�C��!đim��%�Xmվ�dv{��<�W��	-�sK��cy��`�[⋚зlV�{w��0�g#V�^��[ü����-xb�34��λ�����ǐw�?�ށ~+ĉO�	�l1S�Oإ`833q�vH8B�3�n�� ������4�j4'9V=�Z�m�J�&��$M��B�T
���!�xNB(�<�r�Pz���du��N��j�0,�h�K�+k����x�UbB	ڒc��<�� xzz@��)#^|�E�;P��D��v�aI!��㏫b[�l�/a��Gq׆��y�sx��n��Z�ւF�oeR�	��ܗ;�c�tk�͏���Y�aI�d��$�0_�I[W�c��c�U0�G��)0l'���y�0�
����a4d5���y�_���`���+���������ل�/�q��0��P*��>��<'ǂ�7(��r*K>��jL�6��{1�c"�\:/>��?~?�o^��o_��	�p�������/>!Ѩ�8��]��i�g��Y[Q�&�=�P���2��X���8JO8�-��ZQ>�-����Ը06� ��h�DѸ�׸1��� ��p��cV���������� ���T��H¨��]��C!J*��t�:d��"��%��l�,��-T-l��mg��x��U3b������`�3X`8|�5Z�
���sR�R�IH��8����G������ѣ��bU�� �����x�	Ò�8���������|��I��넯1�m?7Ǥ�9�J~a�Jҫ�cy, ,y�Ř�ōz��}��# �E ��o�1��r|�x�Uz>sS�UЋ01��f��0�I�#,k�94|$�E��&,�O�WZ/��C0,^��#`��'0��`��#�1>u���BR��r̒g��M��{�>�>yFe�p�0A����FWa���={gϟƹ�O�җ�a����H/�Dn�,��ʧ ���uL��0S�����K�����V�RIUA�T����Z��a�h�>���&�P3�G�$�͆�0lk�+A�ָ�ۅ0J�.AXG�t6c	Ò���VAx�tXM��OBr�<$Tσ�lAs6a��AZJ������a��0Lؖ"
�T~a����&�z�uKT(�x�u��a�'W/V2��M+����E=͙���v�f|	x>�z���U����H�L�D~�b� [��+%�	�R&�U����V��~h'Ǹb�I��t]!�L���u���b-�1��.���|����#��}S|�b�p��z�׉�X3��ZLFQ-|�X�<7\R����ለ� @s`��m�AG��p�3��!�������bddd����+�����:(Q�L���V7���;�X���0���"�4�81�p�.o���^��x;��|p ;�{[_ۃE��=����)y-X~ǣ蝿�4�q(i��#��`�G����x�ͣ�w냈�υřO�(tN�g_��/���I.<��6lxh=�y��z�U4�4���MM͸�[p';o[��$�5���[z�޾���)�{߽��َ�knó�n��yl���2:�.���[l~�Ud�M'K�|�0�w��0�F�S-'��J��Fu;\�-�XB $�!�s��B�xe_�q�!<G,�d+�ECq������A�O�͹�KfY����zc<a���a�#�ɉ7�F'#nFN.�&L@K{;��kav�M���m�+*�����
g���j� �093����6&Ryz%�W��F]4,F͠bQZ���V`V*�IE�|Y���B%�%�Br,��]*��P�ᜌT�q�o�Vb5��cTL�x|5�h�$,B�U��Z�^<_j;8)ˢ	��`)W+韤<�Ν;U8��6��-q�� ���B^���|$%��h��0M@��Cb.l�U*�_l������x��x�hի��R\RC��M�_�x��m2>V�����i|�ם
�0�Kr�(v�r�%�7�i�s
LjBt�4��Wc�C
f�+��̟�����>�p+�+`����a
P �w�;���D~�U`|M�Cm�g�g�W�S>������k$�K{�b��������~��ģ8���8���t�^�9,��CVR2ۙc=�#�c�O>���BNu��ႶY�i��>��9B�=��*C����4�J� H���ͦ�#i��R҈�I�X�d%�.[��4�%c�3����e#5-�Pl�MB�,z��h�g84�m9J�FH[�6=�	��݊AL�5�5�w�ODc]=
�h�&BG��񾩹e�
��؇��R����@�2��si��#;7R���qB�ĒJ������o(i�xL��7Yb���,�gYxWUU�z~~��I���F���wa��[�x�m���5� �Z��R�g���TB��%aWe��GxH#u�*��,���7�{xH*~�TFhC�������I� axaX*ۍ���sH
���i��nx�΀W�,B�A��?��i�f�){��!@�g�"��K֭Æ-�������p��	��(��!����sgq��i���.+~�Sf#���KQѵ
E��i� �i&�����@Z}�k�#�l2A��ŝpN�������E��ʦ"��K��L��x*���p��"�u1�&,���\?��9����`������e�~�4tiÝ�Ṅa��|L���pk��"&+P�kb	:9s"������
Ã�$��0��Y#��X���K�����a>���u�T���ݑl�#iI�fǑ|�VN6�jxZ9��0:��5��2p��$�o����b�T0s�Nm��Y$�UL)�8,���%�+B�8�`I0�2g��,�>��@����x��@��KR*L�d�p��c�� k�"Fo�ծ��B\|�Z�t���u"fΜ��sb`����S1\]S��_\�� !X/�8�G�B�.)��e�q�wr@����U��W^y۞߉��ÑQ�H��R�"�}jf�e;�����$�[V���j��'�|�o�'�N�=�=�v� G>��C��ĺ����k�س{p��x�ѝpeT������>�}�?�v�;�S����N\A�^/�#<�1�w.�|�#N}|UM5�8<�����d.��'�}�<�}��t�-x�������߇9�cWr2n_�gΟņ�����
�e�o�C2A-�`WE������ba8��'P<�Wa�y�	���0Wa�Q��,搸^��WJ�6^j��v(횯WP,�sC�;$y�֟���@�R�SʔV���R���� (�o�PNFR8":�������	�Q�A('�(���� 8"�F�*�a�;`4�Tn�!LJL"�9�F¨���,�8I�ų+9����->g�*�gX�C��W���+�䘼F�	L�h��wX�%丼F�%�X�I�E�Ã .�xa	�pK�b-6��ZI,��L���4���@xr1b�����*�֭[�����m����J%�D:�N�[|�Ш����x�@����o��at`,����ߜ���
$�sF��Q����A�es��s�2�M�d\o�;����0,�,�1l���b�+�3�Wa�O�vű,���v���7a��˾��ä�ũ����V�l��"�0�Qҳ�v>�	�_�;w��+/<�#－��#Gq��7�v�JT���[1b�=�ع�=\�hꞇQ!V�d�p;�,#S��e��k�Ǿ�j�kRFJ�R##��U蘿O�ڏ�.����8w�"�{g?�|b6mވm�=Ic�%�s��6Y�
oܸk׭FAa�����Q�Yi��ac��^Ú(�}J�գ��S&w�������`�LHP1�9�& ?y�#l�x$e�-�~BL�/��i���";?�F4A=#]�-��<�5������eHO��"\7)CZ����Etbd.Y�Dek���E��We�?��>:~Ol{Eu�nŘ�x�0V�C���`x�l	��RuP��#unϼ$7q/�x��s:�;	q���t��s�-��}����5��y��遟�a\�'P�%װ'��Bbx�T��Tx�M'(���s�g�0�� �ٍ�����ܸ�V��vg�!�~2�Jiz°�c~���8N>z����������O���ᩳ�^1%�����Pܵ��� �}>�Z	�-s��:iͳ�����0���YH��z�7���s��4���Ab� �>)��d���n�ʓ�Բ���n>�|�Z7� <����R3ƫa�a�� !��!���jYL�c�L�+�`��'��[̒h>�D���0�3��I�M ~����%}U�ޚ����0�,��j��e�RDq�M���Fx����^�q�^v�`��n��t��sÓ$�	����R-2�:ZK��*U�pi�*:�Qi�W�X��E:90Ɨ"*�D��r_c/F�� ��d��`��k���'	a��M�`�bͽ����H�̇FG��KF|B*��(,���O>�� ?��8��<�s�N>��N����o��bFhtb	5��́�)�x��]xc����ʫ|�Q�������w?;wB��Y0�U�Y>��?������P�Lz�|$W͂�`l��$�sЊ�G笕����;v��X���X��f9�%N��{ޕ,(�����;�d�F=�-�<p�KQ�2;�:��<����"ڜ�q�ј1{1.|��?v�e{-z�!,������xc�^Է�b��Ÿu��X��V�[�s�o�\�ϙ���t���V�<}�lX���"$&����-�NVl$3��Wa��װAep�p��f�9�)�Z�	�� 1����\�k�4�J��R<]��Sy�����S�/=$WL�<���uy�^mFR����9�%+�aƌ��>�˖���w�E{��Λ��9s�4q"ڧL�-k�`��c6���
��~M&��a�%�<Y�^$��U����2�����L�5��Z��X_�%;�*B���[	���pC -��! ,�a9.[U~9<D�+�r�M�9`	y �
���[r�W&i�
K<��L��F��;-�AA�a/��8��F��f;x뭷��c��Tj�ђ�?%��;�C��j�I���3��n�Ko�o�U�=*G��)��BD��"&�E��!���4�4�K�� ������waX�2I��*�QB2�H�9ka���L�*�x���,w�"���-���!?�zϲH�k�������0,�	OiDς�p��E�Z�����1N���*��:��O�����'������Q��_���z^� O_⸶���_�ݐwU�l�7�^���vİ�kr'S���2Y�&���Y���މ�'>��c?��)�x�<��}xv������3ܿ}�J���6�)9r�3���G�8c?a��[N�7�B`X��pl���Ϭ�n����a�0�$UjZ��H:4�3:�)YH�LW0��T��#��hu�HK�vu��-�f��V�$ny32������"K���	������\��ҥKU��B���<@#�)ܻ~#���*{f�:g�3ʁ�����1����a)�MI؃ ��I��h�ǒ�T��U��u�W�FM��<q�ٛ�8�d�,��%�#�,0�s�&K<��pa�O�r�M�gf?���@�^<w�^�N?��ْ��Y�Ƹ�nܜBv5c��09'8�I�`Xy���>r�&�׆ay�����U�x��Q���;�ξ%H#�4�F6�%�})���E��'�:)a�E�uq?�ۤ���{+��ܸ@I��r��;���Լ������o\�-��`�!u���$+��$���g\�AS�Fb��T"�Ed��FX�us����VHln,�,�<+�Xb$�0\�����)��%�0A�0���K-p֨���w-��~	�|1�5�w/�D3~��i��&r{���[��0rM�Ċ���RGB�|dr�Z��#�4���5�i@������ �/FB����ʙpT��F�����i���v��ӎ��Ipp�;�9�s� �v:�s�8��Ǹ����r������/��:�&�bK�NG NEt�	�%�j�ԧ�}�o��=�|�>�|_}����;l�� ��q�#K��Z0;���u8v�".~���<�+�̋.�ĉ�8{�s��S蘹��f����\ԅ��~�s�h4-B��[��vQֱ�ˡM���P*����ޣGѻx*[�Uz���ơ#�q߃/`붽8}�l~�����w9�<�*V����������9���X��q��U#(ڊ�+�����ȯ(B�&>� �X�۶����ڃ��FL�я�+oǢ%˰t�-X�j%f͛���yHHL�-�n���{�	��� ;/9���C9��С���/�y۫ȩ�E�� !4�"�. �Њ���p��q57,�}�@,�/���"(661�z�(��8�u��N-�s/����X��톯1�P�}%��ҩ�f�]%Ȯ��;7>��������8��8���xs�>,���]8p��7?�$>��/����0g�|mp���0�%T8G�J9&��S\���ڐȉN`87�'�T�x�\	�H���`�a7#-ى�T9����O�V�qr�sӒH�Jz�7ج�I�Dxp�Zlg $K���L8��
�%���J��B��V��ׇL!8A������j��@Mh��w�/)�"���z
?�����~��q�{�j�NNNVyQ?��#5����ز�Q<��q���^y�m���!,[�0���	��
�C���/��Ȭx��8S�`��V�`���0,c\�06�a�t�`X�$�r�M�!�%�!�s	�C�V���JK���^�?�aj~��O�Z y��{�~�2�0,`�����~�����X:o�c^zl���ξ�؃ų *"����/䔔c�Gp��0i�
Ri�pN �&���a.�����W�k^C���^�$1��7<��d�UP�)��p�}c���Z��$�䦡����'���
ڛ�?Ѓ�n���,@&�@�`	!TҧEРs�� � ��pE0&$�cu�p����!,8�A�T%�T�p��ΤD��'S�3����N��~����b\J̰lE�r�Eb�%5�������K���V����IE(�F<?9%�cl-Zih���c���X�\�y*J˫0�o.�X�����'c�,��JU�3�Y���D��҄P9��n�d���C��#}I��V��JP	Ir{��^|q����U0��>�rv�-�}�
���tEKȖ"Rl%<�0�9^7�5 ���ᡴj�ky�^�D?�����Q0<�0�<Ä��NnE@�D�d��&����ٷgO�U1�*������?�'OƧ_\Q9W�f�P0��0�L�pz�R$���w���:dG���|j�	T|=��պs�Zkxy�a	�Ka�9F¯�v���8���s`!�/ELXk9|8�'V!6��@؉�-Ϋ0�k�,ت�|,����*aR}NK�����°;DB���[��r��<�7��n��S)'��N����G�p��E-���ȴ�T��.�Lt��;1������ɰK��|��܍��UH�����Ǖ�U3O}�x*�n>�������`�sv�.v������ip��!�h:��EyS�lDc�-�w�����=��������x�����a<��a�g� V� �.NW�8M͝���A��w���q�@{��iUiP�bϞ� Z��uaI3fv&"��対�Ǆ�s/��i���{��x�����1�w%�&�Uޭ~���n�!�Q3�v+�ؖ�_�.	U�x���8��7x������8p�N���l~�c7�/\�C�?%�rP��@E�d�Vw���~�������`ѪH��57�g�|p�4�����K߿�~�����>��(�{8����˰��G�}�.lx`#֬���#5=��_|�5^��&O�BgW'��B��V��5��2��ݽ����_�M�$,0�6)������T|3B�X�"����J�Px���X`��6�=�s%g�� FI~��
&�%�_G��H�A�5����m=�4u.X�[�ߎ�sb`�<䕔b�����l6�����m����><�أ(��B'�Pb$'Q��3�8љ���|� +5.�.�i�Ȝ�Td$%!5�Ev"��j��":��&� mAUEl��\VR��M�u�f�g����B�t1*�Xb�%�ZH�/��C���[,�-<�6�Ey��{����N����l�#=3q	Nh���dmR۠�P���Q�,�+���Ç��K/a�D�!!
���ʕ+q뭷��kk�܁3z1�k:�{��5E����a�=�0\D���HJq���^���=t��eIo�x�Gx�C��!�0h���p�����A���2vaH�\��<��\B!�8W�x���տ��<����ω ,�b_N�"�ò�`�p���`W�ͽ����|�������MŢ���r�=8���:x;�{	��e����+$e��-;��7��*��,��H�CHJ=�s��PM��(C1n���HJtI�/ok��9��8�q XcE��Ʊ;A�(�X���c�V#`�IY�X�hb#�N}�#<"�O�EhnihdJ)e15
��ek��a1�y�%�>:"��HILb��A��"� _�H�HG2��}�!J��Z<G8Ix���;.r����VPl4�T_�X|	�
R�3�����'�`4�B>�5~��B�1���P�v��29�6����������y9��T���l�& ���݉�A�x%�� p0�Z�
*!2~���]`����9�E���2���љe)�F�N/�!a8m
��5*'�h}�`6�
����v�a8c:<��9�Rl��@X������o���aB���'axT��=Á�0�Xۉk�`��Mj��@7Tt�o�gx�ϟ?�;C��W�����!u�2$�eq��`f%��(�d�a�_Q\�b�7.#�.'/��R*���>�k��5-��� J(5��Q��>�c�&����`X�!֤���30l�V`X�Q<iA�� Zs1�Z�&,lЉ5�p6��#��0���C0<�0<���Z��}�����Z�D���4J�c��<���ȿI�B�������~�ų�� �K��2�w�Fݎ���KltA�s)A�z����\+�s7¸@�lͲ`�r'�^4Ῐ��~�4���|�r�9z��~���x O�܊S�O����+n_����A(�~
�vZБT�4㍷��ɧ��ot'Ϝ�ÛCY5C�� �ÅP�z��6<�w�/��:}x��5��;pnzwlx
���٦�"���.
��\X��T��2N>�V��iT�k	fg��:�}�A|������?&�>�*:�̆+��Pz+��m/�CM�4$e�#��E���яUw<�����㗱����U҈H�Ko�����O�D�	�cp�}k1k�,U����[�Lʆ��DeM�x��$��W��|X����8w�c�e�����/�?��/nCQi!
K�{��򻯱��7���O.$���g��a�VD$�"\�q`�8��A�R�x ���R�jhq\�ܙ��-R�Q���j��x0$�/'_��
�#Ȟ� c*"ͩ3�̈���w ��q����D8'?��0���B0AP+Y#v�X'<�#��$N���	�Y���B�Ӆx�N�)���NIAzb"2S��ۭ]3�V�piL$:�PUY�-۪р��l�����IZ���$�p��;���\r!��7�����ŒY"�fQ,)�sB�X^�BI')��`�NȨ��CN^'h�:&�����a������c�/��/*Vx���2�	�j%�L�r�W��1��hb�Y��$P�c�o8<�-�f��T
Þ�a�!�a�|:<LZ�R����M
���0�qH*?�K>^	�����s`xx��h(4B�����i��Sfѐ>v�N�ǼYs1������^�Co���_����k�?q}���摰�����x��E��M��ϘD��o/"��Ç�V�U�ʔF��s��'X�Z��}�G}b���G���Qc0�sa7��3�����ia��E��S���%({(6�Im@)�,�>V��}�ƞ �x��Mz���}/U��(+.GeY%&NhW�]ŉ�������@\H�5��]�G������E	U}G
�H�Q(���TJ���4e�z�����׿ň��`�Xo�IA��4#&!O݈H�BǷ������2�J���B9�͋�R���X��1U�M�2fJ6��-&�GX�ctPR��p\�χoR="��
�
�=�C0,�$T̰x�	��Y��ʜ��0����U�p׃���[������	_8�ӧ>������Y˯�pa8�}9�ږ�"�Jص4,$/����V�P��Ih�b�t��jnk$6x)!o	@	|�x��RK!�����PC�	��?���Dp��I��U=�'0l�a�9��P�dp��jќ�c�8������23�:�]��r��°�g�Saa�N+/u�,Z�]��d#�\$;�X�������߃�� �c��g#m"	hZ�Ԗ%HkY���$7/Aj+߶[�޶
�S�!�k��"&w"0u2���a5�a��Jw����C�r�Fzv2��b�0e)�$A��x�����w�g�L<��8q�>��2�|�]�j#L��,$$��dMF�ƌҊ:<��3
|��X���^�_}�Sl��-���i��]���cr �`��%+����p����C���W�����H�|k6<�ƩK�X2I�����m�|.��&�[W���?6���iH��KF-J[����'������;p��'���-�ȫ�і��˰ｓ���NUMP��_�Ɖ�H˫�9!�n���_��W ��a�x�Xs��8��2q<�ǡ�P\[_������S��э),�gr.��D�n�&��	4��n&߉�}��Ӄu���#�me4f���C����f��3z�ð,�kq�pb�Z�2Fp�u{|ݷ��X�@qP"�W-|�wg� �Eq���󮓄���"PK&�D�)e0�W��X �+������D~��4�\���HN���Se�0s��5M���Eg:)�l�Vg�Nˉ�ivF&a� ��B�ق�I��,�>�`,��ܬL����HE�5;+��*q:aY�?�f�ns��$K�DAW��I����v�`�j&	n��#'�/l&D�pb�xr�3M����gcR�T��q"�W�uz#4C0����������H��ܹsQYY��yq��sRR2����%5hH�>y���H��� X�w����W���I�Ν /{�
��(Waqu���a�����AC0����0,)����]`8�0����y�����㰔z�\|N�����g�1y*&TWa����؂���ݻq��i�8|��	5^㑒��7���Cg>AQc'�y\(|�I*�ר�D�Q&Rq��|҉4�����>^�L/�{	l���!P�Drn9j9f�5���99�HKw����jc�u9 �����g88$�SY0�b�=���U[����(�K�#V;i��#59�%e(a�.,,D%��x�m���r��u
�u�\I��K0,a�3,�$$TB���V�q���aLc����'������MMG���h�
gZl��Ȫ�sv=|̹�0�b,����|���B'���dK����5�#�Or1���]n��fC	n�cY'�%n���o#3�m��T�opxz�d��:u�H����9��ݹ])��vx-f�O`X�	gO�
�?��k@<<�gS�� S�ð��aI�欚��+p���v���֞�K��卮�&q��)�!K\��b��2�VLBz}?�[!��2�0l%���(I�3�A��ؐ�����f���Hl^����H�D�kJ� 
�"�f&�
:�Ȗ�=�mY�D	�(�}�L	�	�Rt�vܶ"��ڋN����Er�lU�T�"�Z�����>$T�ZB��Q	U�$��'�U9��݃��9�k�O(�?'���,�;$X����d��+��	rTs�P1�h����{j�#s�*$�x�4qv�Ŀ�\=6�������s�>"����;΁�d;�L��̤%9��]2�л� �� �N��c*������/�w*�Cl�tD�O��x��9�m۷��݋�y {�ݍg�?�E+g#>9��,|(�ٚ�)����Uu������a��سg�?�G�|vW*���1�	���
�+Qz�J�6�o��A,[�Onق#~�O/��6!��iM��� �z�Е��(�:�=���^C9�2^��~�MA�9����������`܎)s����Ǳc��Xp�Z�7�{`)^�=�Y%���6l�<�uJ�mME�Թx��i��7LE�9Vދo~|r�L鞎 ??��	Н���%�T!3��ߡ�0\B�!�1i��)'�5ɡ����Y�0p��k���\���7v�ҷ_�W�AN� |MgU�0��E""��r{��C	��[Vb���6 K@����4p"�;�
�E�>���^���S�(��T���e���=��e�MDj��y�l��x�l~�%<�X~�Xy�Z��a�w�N���v����z�y�[�z��a�hc�%�t��4����
��[�b��Q�s��۰�A����MM�ߑ��7��-�&���B#�	���J�9ٙ�*�8�nQq�K��D��x�#q�v+�נS����f!�b9�
+�-'e)M 0�ܕ�������NZ��G���_���4��d-�zd\��Oo݊4��F#lv�g���＋w�<���&�w`6�g#6lzѐ�Y�ƌ*���y��ymja(��؂Nx�=�E�!,y�Upk��@y�ax(L"�Z�r8�٪�h`7r�-�Ǭ��Z��%�d,5��R����D�NE4��0�1�_��ⅇ W�	P�-��?��0L�{ ���?[`�6*0�|5N�?>�)fNꆆF�>4�N*��ۚ0�{�{����#�!9=����9���v�+a8Ș_}*���4�K��A�z"獼�e��vb2��#��x�Gp\�&�c��k�A�?p�8�w�އM���.<��ly�ܳ~-zz�q�-Kq����z�m(--F��.���Tj�CXb�U|���$D�� 80H���(ww��/Re.�A�Jk,ƞdX�ج*�Dv^��fdg)� ���!�]�#!�!�k�*}���?~��_�ju3zf ��@�\�W�NJ�'� ^�t	f��`�N̞��_|�^}����cO?���Vcź��5o5��
pCh<��faaxa؃0<NS��1�c� r��o��č�4Lf����E�b�6�1�A*=ʂ:���%Ps_
��sl�����xUg-#���m�8*T�D�T2�a��f�*fX`�������pV<sf�ga�X46K��]�`������:��9-�?��"��B�n~�n�N��ffN@hf+a��V�Ě�6����R�$Ο9��$NK�0a�¹�HF�2���
�
����E��?���N*��0��C
�S�i�HS0�L�x�-u��z��k�c"y�-9F�Y@���hZ=���2'ACkו3�-p:+a���w���[ѷ|�Z"Ab�ea��ζ-Cta�Q��W��*D����f]�ᒙ��E3U\����>d�����p�H�J�t$�j�`�ꃕ0�%.ПB9j��P���f&\�e{U?|���TLQ�ܾ&��2;T&��ɷ!�c%4��]:Ce��	��������i��"�-�v°�r>��`�:M`�t���K"�p."���K7W/�{.Q0U� ��sS�ߒ ��녁2�Dl�Th2�T1��چ����Q��._��W��^����Lqr0�q�OGTL<$�:+��lz�!���؏3��c۶gP���5a:;|"�7$����XS_oB{[6m| �}7^x�	���t�r$%g#3����
Y�S_H��@Hf��g�T��F�J"h����DTb#��t&͹�?����;����(jnǖw�إ���ۇ�j�&<�������!L�]���{��o:���e�����[^ĉ+��6]U��_|.:r��s����Tg2\ɰ�0�u:4��I��r�
O�FSB �#�%C�s"FkCd�	~�� k&�Jg3�k�4��� .~�5��>�Ҏ��7"�0欥�lK�����&A�=I-���������
~e�GX*۞,��� B퐮�s
& �H���}�8I� Ǧ�͙Ȯ�Ʀ���k�/`��'�֑����ر�^{���x���>�5��Ͽ���x�8B£a�%Pq�Z찘����0��`5��@l����F���T�1B�H�=��i�Ve���ab��u*U�V2E�@r��~��u-�����C��_��K�Y-�#(�$Փ�N�}���#G�۸��]��\� -������E�eT�{`�}|'�]��w�gi\P��x�@s;�>��>���nĤV#&C�:�p4���3,��$fx<��\1�a�ð� K�a�� ��A�V�_�aa�Xp�epda�h����Aa7�<��{4��B<~���l�KZ0G=�3��ݯ<��?<�YSz��@��Q��
��f���C8A�/ c=|0������g��/"�j"�ul8������LD'V�C�15�Ee
��R��F���ѐI��7a�ל���K�؎}x���8x�<Dދg�}/��v�y��yO?��ݵ����m�c|����={�m;V��e��*�g�C,���*!�a�#���_�	��lꮊ���D��Ѡ�8b�`��JVy,�7$dB�}����������J������9T��,�0N��P�{VQ�,ƂE���O)s�[���pߦ����M��4&"�Nxh��/�x����*���"�J&/��9�!�`ٟ�Y�1��;�X�ђ2��:"�7k��"$��W\�@�����f���zB��~�lG�3�+�Ɔ`X�.P0��a?°��0�ָl��!�=��'X��3ݭ�{*��t�
O�W�T�N����&�p9��0����[oŝ��m���7���G'_����:�#��W�s���S/�����(�yJ7,zl&��}���.��j.�E�pT�A}��܍���3ofκ��ne���~{�_����Df�<�6��k8G����a�Q�5��L��e}��aI�_>��|9�-���X�����gE�J�e-����r5-@�,�����$5�S��'U��u����)�5��D��{Qر
9��x���ט��̇C��m�Ep�.F�,D$�'����e9�sF#!��Od^"��)��H��,߼����V�GxAx6�J	}0���s��;M�#L�`J�3��˰�ѭ*c·����"ڻZ�;���/b4����'�98�;�p���[W���c���E|��E<��V�VT�u�tL�9�q���zG:���h#�2��ă���o���'���m
~F��@rF	&�,C|N�D&��W�iEx��.AB�*�y���^���X0 �ޏmo��$������[w�vj?�����#�~��K��_Ǝ_�#�x�],�k�|�}#��;�9���G.s��W��f3,Y���Jƴw�2��G�����ؿ�}���=���m���u<��6ܷ�Qܿ�Y<�䫘1�8h�EkK�5�F%����>�8~�ܹ~#�}�l��<�'^x�8���{�7>���N\��8Nn���-n�p=��zI��;	�r�M� �H�É���Ã�|�ý�?��K�0��°h�Ÿ�ͬ�XB��5yP8q 	%-H����	Ȭn�q�MME\V'��[��?�4V߽���1F�F��2p��s���_Bm�&��A�Ͱ�-�b)�zf��[M'QJ�y��@<\<&p�^w����$,�?}ޭ�aX&g\��z�J��sC��8((����U፛n�	ӧOǛ���/�H��v���!$B���RT�LG]s?*�{�3{f/�M�s�,����\Ԅ�VZ�1N��k^�`�P�E��/!�ϰ�z?W�J�f��!K����_�2��@Qάk�����:����	�W�؅/��g?b���xh�Z�\��W,­w�֭�ʵ<��.�ߴ<�$^����s0ʩ���6�φ�.�\D���C(����߆$�&ߒ�(:]Rl� (��J��@K���1k��xx�Sظ�A�왎��l���$[�1�U5娫���e��䓏��7����c��+��f�g���4k�4��})b����.0''G���Kֲ�Iᥚjd���n��ab��{X	����[���k��I��'1D�&L@Ii)LRЉ.�#�-k����߇��F�蛉��=��#-�e%�g�ģO=�}�3C�\_C:�YT<9f{�1^A0����f<a؃�:��H��؛$�A�f����ޛt���h�A �7�+�e��R�EA���K��/}"��4����$�$\�a�����#$��y��ϝNx�%��o�s��_���O
���� ���p�B$�paO@�n.d�H�E����xL
g�I
���]�<^=�
��8�ɏ��?�������p����Hh�u�K�2]|a�|&t�-��]4�q���H�F$��0\; 'Av�@��"����S�.߯q6\5ZA(�����k��R?�m��nS�Y����R�
bh�Q�}+�W�����!��i��霃��.���湾�J=+�)l�������7[&���R� Qy��%sk�fѐ����*�"�Sڏ���0�O��͖5��.8iY����	H��D�B�w=���_Ň'O���EZN2�'7���#>>��Z3�tI��5 5p�|��8��^��Xw�����.�@i};�#M���)HH���eDx`�e�|�>=y��1� �c�@�1#��ҨB`�r}����%���9�v���f"4qjz��������b��ݘK�M&���L��{�`�#۰xÓ�}�v���6Pw>����<�7��9Qm�܍��m���>��ٟ���[�����<��K���?�����[���p��8t��~�5>��n��;�+A,���ں����� �㓯���_}��_~��_|���|c� ?���8��X��H'�D:i�Ѡ�ph��3&�\��x8�7��b$�J�Z݄0�
�ҸO�{a8���L������CA�9�" ���1�`��.�U
]Z	��4
�m�W� �����C�>�x���_ʱ�h\��h��d��$^a�Qy��-z�b��*e]M�h�,+�%&X-n����H�)��`x���_��0,�+�Lʲ/��V�x�d��T��TjR~V�ˢ;�aɋ��m*��Ƒ#�������>N�>Ai��(3<��sT�j���qAx��lHQ�$"�%N(���}�I�MVa�6^G�
��I����c]'��0���U���I$����`X�W���W�P��y��i���,�G�����?�ۏ?ǥq�����c�7_���ǅ���o���?���;���G<�J�`�_<b��̓�>Q4x��d#�^I �<�y+:�Y��)j_<ã��8����q5ʔ [|2�X�q���Ap%�!9�_���?�*�(>ޡJ0���p1R�4PERny8ki���u�����SUq�Y;��/��d}��V�YYl��*�Wb{e���@�����S�������h8Ο?_�����N��%l��Ob�G����U��/�_e��/,P�f8e�Ť 90$��y�+�ڒ���fT�I��
�+��I`��ɾ8N��Ⱥ�>��>�15:{�8��%r�N����x'�a��ޮ	�?nG�1�P���ոQW�bK�[M!���<�p���l���O��E�x�_��>B矗�(�� �<�9h�k�OaX�$a�INlBP��I\��?�Gç��0�5axϻnN�ð[F�iL~'r:��q�����[O����ċ;���/��}�ƙ�����F2��Rԍ؂nhK{	�K8HO!��ÚG@�R�x쥓�Dh�s0�P����ִ�ȁ&���&$u�IYrZ�M���`"\�S�VӋ�����n��ڠ�s�����B!��Z���yh�Z����(�����~d7�FJ� ��v6xN^NZ��Jo�F�9!�`�1�b'�tH�*��"�N�=��i�ʜBP쇅��/#�@<(!X[ң�+�sn왝pdv .c"2'� U����{|�<�� ��{�~XDj�����,@�&��>-v�6�K-V(*������{^�+;_���WB�E���L��P-�1&�	�|��1��>���އ93zI0�! T��<#������&�^�$[Y��K0�����=͜�Ó'!"��	�Rč0��7�
k%�H� 0prO,Ct�x:ym��Z�^�P~N@��~�A8���f��L$�u��@TZ;lE���7���f/݀�?��o��E���.Z&u���-}��>�vd�/h����0��V�gv-f�X�u?���?���l�v�ܷ��oƪ��-�����d�#(i@\a�iT�[	>�C.��� �<�A�8�3'�Z����^,�8���H�X`xH���R���J�W"*X��'� N����S�����w���j��4NV!�,�Vw����q� �*FN
��N��#(���(F[
�FZ�D�mN�&4z8�V��%v�J�Y,H$\
GEF��f�x��bYd#yL����$^-T�*�8K�`)+k2JI�ñ�Y��T��7*JEpR�����0�q4?G��W�Wn�A(�x�eR�ϒ}�`�! ���3&^2���駟�s/<�<_������L��Yi�iph+`M�s�$�iJ0&(�\�� ��0[�J��*�7�{Ѐ���P0�a/&�KU��7��H�X?s��°�0@j8k	�N�R�����\~�=����@q�-ؼ� >:��ίq��'8y�c|x�,�9�/_��>�k�籏�����k6����y�Lh��㿯���"�Y*�AP�j��)�c�f���"I��k)��,�%s�K�H�P��1��FB��741l��Hp�PV^���#_?o��P8�l���h�O���C�U�4Y8�aw\���h�J�>iDnn�2���PL�MOOW��1�c;:P__���Z�MhCVv�����{���R�<��F��%J9g�=bh
K�)�<�����G�jMb�{Ӎ
�%�X�:53C�'%��B��|���������'>�N��t-y�������Q���cAx�N�� ��I��S�h�:A$*"z�3���˘�V�4��4��A�47(8�QW������������V�D��x�7���&[ �a0�7�9n� {d��9@��W�����?.�A	+@տ��ؽxN�=38&°����i�ҁQ�fx&6+㜖Z;��s/6lz����'����I���~���ax6%�4%��T����q��]X��c�똊��bU	͕���	�ز�-,�k+'\�R�4�9h���aX��p�5��йaX
����$h�B�.��m��F�L@jy�*���܇)�FK�J$�L���]�҇Y+7b����M֧ 6.G.镨j�����(����i(��En�ėt��e˅����Q�0�[��a�`=����MFb�0�ewJ+�o����߫��Ie	In�*I����P� 3a�:D�	T��p]."R�/�Wmf�gx��xiכxk�~lzlm���G=�v�=�����5V���~(�j+���Oc�O�U���{ש�Z�%#��x��X�s����@�D,Ay^o?��܅�mK�"<(���������xD�E'�#�Rc�D���12L�S`-�B}�������b�	�3	�݈���4X��p5I�A��l2�����D�$�˥�t��SR�@W8��b��z��ܝ�� i�Ҽ��E�%	��	e��3�;^�T0�q�:���`�>	~�bD(�y�`�jE�@��(�c���Z@���X�m����8�	�8�E'AKh�+��ϭ㤗�IOn]W+���T>jۄ�M"�:kL�&��;������/(�:���`�R���mN�gV!�FbF�|�r�ԭ�p��ea�&�s�KE�.��1m`)�u%<8)GA+`�,RB9�:Iפ#��0p+2�b3�x]�Rݐ���#$<RY�"zp������&�A����#���h�^�I؅�`�$�@3�(�	��y�)��b#�yٗs�%[������[�U&��I����Qe�����447�"6���H/��@�)��Y�p[I��$�s����c.�@��������Z��
��YG��a0\�B��0l�q��(c�?���w�aw��$�xs�͙���>���`��9��=Sz桦s*2�Z��҉�I=(�ԇ�)�잃�isQ޽�mK`��6k*e�ׄq�rxP�&�����Q� ������[��?:&#�pS�	�l��$"3�UU5*�3����v�����r.�A`��3>��P{�#�d0�mt�dh1�n��������Q���#1\�ھ�ա>#%��%�~���1)�CS���bL�sr�<'F�x�e��_�J���7�}Ş�g�� �J̰�-.�!*��
J�Q�y���%(()Ge}2+aM)�����{�s�b��H������������%��lQ��k��I����)�!�d�P��������2ͭ�.x$�a��7hKĄa�x�����]`8(�0���0<n��a�<�g��T�3�@<�Wax��p��aXe������}w�[�-��!�qaxս�q��M�㮻U�s�0,%��g��<�	"�_L�v���AtpBK��|�ۗ�;aX23�D|�d���k�]�����#)�)9yH�)�+%	i�h蘅�)��V#�
=0���P�׷.BL�Oa8"��@3	��a�r���-�|�K<�Ò~*�F-L������oE~c���0v�?���~��^��{Ga}�{�W��K�aβu�% 46��,��KP^��؆��jd��!9�W!�)�����eJEp"A�YD/�5_�pZ��r���JD%U#:�!N��D>���dEq�$���V9�-�,%%e*�wl6�+����LA��w�!	3:&�����^}v�����A�m4�9H�s �G�3���$L�c�Nz?���Fx�|`�Z-�p%�����T��Z�!X�խp�,�N�ƫϿ�����Y��W7�� (̈pB�&���=4�H�Ax��P2��&�	���0�̂�x>!v\��!��6���ZŶP:��;���̈́����I�V��V�g�\��!NR�U�A\�>?��y��m4,G��Zԃ(B�3"
j��t��kwF�Nh�3	��	������Ø�k.��4B�-�@l����פA��E�Ɇ6.��|��
��@G�֧T�Ȝ��-��(e۬T
#���@�d�� jD(ˢ�`Bia5<��0�� �����`h!�b�FDf��&rۆ�	�U)h�w:R��6ڈ��6�qP��#@��Q�������|�{��5� +�͍���DEi9J�J������xdef��� �))jb���S�����s�=:Ԃ���4�('��ovn.*�*QV^���4噪�(�qW���<�\	�r��ɨ��Ty�s��T���L�de +#Ņ���y�8��%�w�^���V_��+�2$�x����RuL��I{ʔ)���~Į]/���
�F�d�
AN^��H�;���� N�6������� C�4��O��42��T��~�g>�c��c�5.��p��e�IeA���H~�x�����,LBҊ]b7�_�m�=a؇�yP~/�
�#�`2�8v�k��\�6ى�v�29��!")��"X���9���~\�@��~�ۈ�)�ɝA&"��	e5I���ZCU�c���һ=��nm�67E��ג���X��V<��[xs�{���1�A�n�jܺj)|p�>���q+�L�ļ���nݝ�;w6�\>�8�r�}WD����U��,�o��ڋ���`8#-�}�@��1(�]���b4�!������p�󤰍�@K���4�$�,R���IݝijnViق9O�,q�R����Om}������� ��S�lű��p��i���<�u;�oy�W�ߜ�1�tu�+�ƾ��1�2����}i�$����=���$�Ne{��@Yଙ�����%�d�D ��+�7�����\�#ٷ$�Z� �°o>!2�`9���"&�^�^���0���7x��{fJv�iM9��*��x�W�s/6nތ;�}c7a��y;r\�e�O��! ���_~��J>�0�\݅�~$O�S�uC���p�K�8%�pmLS�6a�yqv>��6m�����p�:̿�V�_�
��[��)<7���:��̀��f��q-�]
�=	������0/�]9 c��"U��f�VAk�T���#h��sn+�y�(k�Ƨ_��+��'.��������ըl��wl�����=�1�6�](*���Z���N�5v ��I9���%�_�@��I��FTbUJ�-C�^NMr%bS���&�U"�^�pZ��{9b	&6�H�:�)TR9$=RB*㬆�U��
�6~������3���X�wL�'�.+޿������p��F#�,��$�f!.ޥ�J͙ݏ���w��O/����֨����T�6�AC��� ��Boq ,�]�s��xw�n\:}f������
Dp�����Q� '`k!UtUA	�����̉���pR&�V�s�r$O&�h�f�P�#�y\�4$�� �@l,���3`.놡�����u��$�o-����pT͇����x6tE�W�Gb�5�7>2���P�8��6�,3�f��z�hO#��Ni��E&���U#���U4���f%?o>,�ň�.G\V尦����%x��YH����K��@�Ĉ�S�����*�AY2=Dr`�NoBI v�7��a7��@a�S�T>[�&��%7�Ƙ<���#�~!�I��q��-C��Q4$�*����x��}Y]n5
#F����UE7�	�*m'\�,er���Y��e�L������J�/1��dI�?��G�iJ���	mN��YrJXBppH F�|#�[��b���/��j"*��^P�ұ	K&
��*F��r��^�yo�S�*o��	��	]�%p�M7�m�p��i��e㷿�5B�O��v�{p�!�4�٥��U"�x��g�sd!��V�5z�5�A��ϒoS��E�Kc�ז�UxAb�+{T9ퟃa)+0l&���*���awэ_Z@�G�2��׀xxJ3��r���{��k�t=�^��ex����A��ѥ�0T�!�Фe_]y�S8v�k|x�s<��uTM�	mz!��2�\K!眒6�0�L!lM��b|�;�需��>x��0�T�є�����mT.~���/OKn��įC�4D��s�}x�s��+���ķ���O.�Ǿ=o������E���M��޽�	�����`��{8�s�
�W:tD��,e	KX����P$
�rQZR��C������)}Z$�R�C���V$�H>OΕ�c�iy�P�e	���x�	�v�m*]��U��#n���T
��yfϝ�i=3PS_�����k�aŪ�1{�2��_��_އO��ĊN�d6�w�M��v��8�����j��ͦ�����X���Z���a|�DxeLVq�*�C�Lq?�2��J L# �����Q0��s߯B��-a�@�Nk'_����ф�1��`8�����!�c�?cc���a�'!�?���t��o¢a0������a8�*Oª����M���^��=8K>����}�;�5��Гr������y��*ϰ�z��2�Ī�Hn@a8�})�[�(O����#L�|���[ݯnثz	!3`(�]~+�m؊���~��{\������?��/\����G�[��FB��h�f �i>b���+N�<Z�eK,#w*�#|�*`('W��!�<���� ���Ox�#xZr۠O�Bk�2|�la����ؑ=I�ݏʺF�V����;q��W���#س��}�UC��7���a��w���q��I;{{�#�>�{}Y|�W�!=�I>3�0�N&��]��'L�d5q�6��Q�!K|slr=ՠ��D�,���9��-�e�ag�9+e�F�6��5ZU��j3�f5�s��X��S;���n�N��[�I�T:�ɄF=�J,^4���ĝkVb�:K-\�I(������5 �`F�Ψ
,��'`���q@��O/�I���Ƒ
�#5E'����8!ۊ���#�"�$���VȂBk�
h�@W��@���i*뇫v&2Zf�YՅ��nd4���ul���L�TMAn�Ld��%L��~z�b���Z��Z>��.�Q��uɍ��� 9���,����E�*�h$����ȁ�>��$� #"!�FL鲘,�\!i���Z02(
c�b���7��P��U��Ȃ���#�uӡˬ��-��˔Bx��ZR�x	���
"�q:š�p�^�?/wH�
��qJ�ː-�[b��p*2�Q��VD�!*��9���6��P5~��}ih[�	�qH,���������ｇ9K�����N�d�E,FM�---�1�c'a����cf�*�*mW�B�]�1w�<��t¬�.�ԉ8�����o�mme���A	��U�g�4��d!:2\Aq��^̘6v�YU�k���T��T�F|���*R&d�L���+��	\B#&M���<���L<��V�9u�ߥ	7������-��H�G����Ht\*��	���"Қ�QQ�(3�S1���0�O���i�����=9���p���&cy4���X���0L�Y�30(0̉�߆ᙄa��6Ä�\I36\h���z���há���c�e������I�\���^��MGh6����ٜ�.�z�J/�ُ��Ͽ���AT"�s
��	�y�S�2���N�O��T��p���S�����N�%�! ��I�������k�9��I*�Ktb1�	h��Ò�������䠹�
�٦'����[p�����w��U�U�^�H�*���ɾ�\���(JeoQq��W�33�ʹ�0d���Ű�x|��X��@��� ��,�] �s2!ƨHR�IEOO&L���(;��d��{U�[������ܹs
�ٴ�����p9�?��މ��D8K�c+�!_�0/�y%��O�f��A��R�ɂ�Q��o�wZ+��Y�	�݄�}��J��ы� �U���*v��1�Y����b���_i��y����un�иa8�0B�&�%�ι��	�C �t=����A�_K��7�T:�p�Oa�f��8ι��!��L��uw�͛�n�z���ޫ0|��	�=�7�a���/�V0|��/���W��O� p(^���!�K� ��6U�V0|�g�{G6u�^>�>�^^8p+چ�=������^���wb�[p�o���`,���{��h�� �����R��J�°�v6!x ��Y0T����X3��lZfm�|���+�Z�Pk.Z{�óW���`#&�g≭����3*��́>��k�|����[�^�B}���,._�ȡ�w�#~�?p������p��y|���oã��eG����j(���c	��1��A��j�W��E8�����T���6��8�
0"�R�H{���Dh	�R��l�r �"ޡGei!�*�PZ��11��x\o�q����/1�'��5�.GiI��QT����`dUb3ƨG8&J��cd���PY^��˖b�-�����E# (�����	�ѦcTD�h�B��$�n�
���B8!K%��v9b��AW���%�g{��`SkC�W���3���#����4-��H�iDVQҋ��V>I����"�i���j��Xz�3��NEgIGd�Z�T׳H�09��OD`��0b@�)������H�#��������׷ ����Rd�� 1�q�;Kb�4X���kV5�	�ڌ���CJ�r��B�;\�R��sר�a�l�dQX�,t�e�ҵ�`�̭@���FDe6#:���ٔ�12Y���@�*E���m���$��G����q��׉Kp��/q�q����G���2��رCA�݆���GW�T���a�}���w�c�ΗUv��w�E#t/N�>���UVUᩧ�Ƒ�G�}�vTT�aΜYػwң4�V�l�}���!�����5��3���Wv���#ذ������g���ӧ���@�� ���j�\�x1���xγj~饗��P���މ];w����hT$��K�CA~��(}x��v�����5�F%���$����><��w�GJa���a����%rl����1�x�=<|�m݅j}~QID��FsdF�c��g�w�k�0|��^�_)�C��K`8��
̝y�~�"�r���
���@��^/�*qWA�o� �����TD�tBK��t�#���c�����`���q��E<	[v���4�i��W!�}*8��K����Hcd�=��SeLFp�$��|M'��I� J���>�\����ט@���Fo������8j�C������XM���h�:����6*%�ǳ��r��c"�~D5��#"d_�ʝ��"n�v��� a� ��F�q*�D��c�� ��F�WY`XB%����eq�x�e!�<'1�R�N�LH��3#^fky����X0��̨hƎ�H���1:ԌQ�	��Tk$~�;��Y��;h�4a��7��0B���IL��TfLm�O�dx�N�G�XV/���Wa8]�	���<>�K���B���2�0��༖*0<�0<A��ބ�1��
���in%O�wa8o��7�
��Ix��b�ݺ��^��1_�a�c�i���j�X°���5H����;�)��]�7��=n>B>6ÿTt�/��! �-� �7�7��p�<>�x��Q|F~y�~TM!�NQ0��>��3�@y\����a7��O=���;��i���a���*����i+�eGA��aZMw��mx��X���*64$�6�'�7��-�
��r���+�p�>�aW�,��	�z����d��G���;~)͜��(	]1Ʉ{�;��Ɓcx�W�6����o]�S��b�����S�sB� �� 6?8��#o�[�_ťO����_~}���+\��c�������z�s����a��F�!�NhJ�����ua��! �$VJ`��0\�hj����E��r�b�Њjh��,D�+U���aK,�6-��h�'���AФ��լ��-Ղ���	� �N�.	�-��|�E7��Lp9m�s����e���k" t��`��b�:D�`�A��rB���ǻ�؀��(���>z�v�_|̸9"��A6����"d��w�Dm���KS��Y>��%H��~N+l��蜿�<�2{�]<��n���X��S��x�z�ë{��7�b�C;1��n$��"�Rۮ���l�wnڅ��{�Ƌ;v�����>~/�ځ^މ�lFQE#t�dX3��@���-��/��w��[�c�G��{�M�ۇO���y��y���+�FQ2	��t^��"�J*r�]l�l�Ф�A �&���?��
I#����J�Mᦫ �`�
� ��sE���A4�T����cJ�!��%Uȭ�C󴩘�b�e;����2�j�j!I�wJ�X�%ee��������*�$�_v�
���M���nU�UJ��z���]L��@4ۛ�"=w�<�,Y�&P���$@?Gx�6u*�rrp۪U
bWrsr�Uz�]�v�_D}}ī��ǁp�]w�P	�� �$.1�.�G}��IH�W��%/��1cU����p�Ѡ�w�����gj�8��e������9�V��?�3�C�ٷ����VN�#g���Q�:��g�Бs���Y��� �?|��:��i��I��� ����8���E6��6B�H�!�ptF�h�N��0�K8 v�O`x��x(��*��?���{d�@H�dD�O&�!4�������ݘ>� 3,�s����o��}g>�c�?�};��Χ`��%��0X`؟0�Oh�'d�=ā|^�8,k2�r�`<�j,���)ަl���k�����^����SR�#BJ�!�	��eX^�a�F��0��AD:H(1B]c4�H�X��(�)-Jr��4H����|<�y�y~�}��\�Ru`O(c��mG�etN?�
�,���h3&[��#������^!f[���'�1���1	����)Bax� &�S_��D�	C ��.���rx��H�e�]��X�O2s�_��^��˯�����
�q "��c��-��t�_T8Q�I���{e��s�K��^ڏS0"�+J���f3`u��O]GM�^^����&�q(/�(S�v_$R�Z5�26�����2�э��� �]� b��U�%େ�a�8�ٞ	����:����,q)Y<2<����"��l�| ���](�&�#{��ENp�W�T��tg����s����C=��pS��u1���+L2��`M�x� �l����B�Iz@�k�1�)��X�̽��Q,�(L!R��O%��X#�0��V���<�7�tl���A���ia5���YurL��heE����X�q����U8lߒ{����zK\�]����������-���a��լ7��b�.�~�h���h>��:?��S|wC�~} &8�cݎw��$��C�y�'q���/~�0<wvk��D��Z��v{D+�~�~�V�����-Y���Ĭ��NƱux�����$���B���v����]s4��4�]����+���涊شC`���R�F����S��f`CVOԄ1ob��3I��~�u��H��W��a)�@֭��'Y"�,��	�5qT�Y�-���>l�"9D��0Y17���:8�(�ʙ��{�{w�#%+G�u(�V������ʜC�4t��CL�E�Q�K�b�C�gE�_m�ɶL�����6�Q�vTC�"�8<@�����e�v�(��q��q�>ٖ�u��꼼��|�9۹��J��#Ng�j4f~V8�p�9^�8E��w^QD��y��96=�*[�8�iZ���������aS�#����~�T�H���y\�^u�q��G^qZ���W��:��C��O��c*���R!��q��9��s��s0uXb��XܟW5dke�� Xb
���>��[���F!�!��l�̄��kؐ��Go���)L�O	U��9�n���xTe���B.B�E�2�9B!Lj7ĩV0m>���d��~���_t�\/����a��:����/�Iw�9m��
u���݇<�wT��ތ�T��]�2�;�E_:�Q8/H��:��OP�k?�]��cc�_�)�m��#�Gv瀬����M��F�=�>��.'de�3TU"�V9 0)VI~�m}�\/g4-���gv�r�:P��f~�� ިvH�C����J�OI�_���
�����Yn-���k���+c��?����@����Oea�ea-'�;�Hz?Hk� 7���R\f�c���<u{�"p+�yw���4\�^�_<�m��u�"�!ר�����~'/^z��(yA�E#���s��?�W��Ka0$��e���\UԁY��"�:W`�zw|�)o��{q�nq/5��&
�]��w-5�^Y�&�A
e�-�U�-��'x��V���-'�\�ϛ��wʑ�3����T��Z��ֶFƴ60AVG��S'�t� �7�fNcHg�� ����/+ uG��98��a�ăT߃�zh�:�^�(lU�LC�xp�F\D��ID�ב�<5�1�#-��e7�On�P�Hm��m^�Ë��iaI�y��o�:��UDZ�ȥ�<5<x�*	�[���4�:1���?��$�]�)��ܓi�*y�N�g�r	Х��C+����*��w�vڔ�>#Z�v������Kz�DL��n������̀0�=߁��x�Yg@�2j�����}k�Ɓ�S���!�T��Ѷ"-�)���`|��׎:�=^��=(T�?���@�q`Z�����G�'k��f�$��V"b���o�����tI갞-� Ġ�)�("TJb����^&�|�yԶ�������SA�Ό�u����a�B�K7����\5e���o��~����t�W=L5Ă���\�U��p�&�S������>�W/({om�~V�p��?�4�S��q��~6	��8U&�Ix�o0>�ϛ���K�yy�z}~�",1~<��\�4׶/�v��e��0u�1e�<��0>����b˭I�U���HF	0)X�Պ��V����v!�eKZbA�r�`N���*[�-[��1�}*@���t8�[	X¥d�E_�xI�b�Vs�^�䈌��~�F�Z֦���1Wf&�϶�sry͛��V�hʯh�}nO#eA{�1��OŨ����e�!{ؐR�,+DO���:6�Bݗ�̪G��7]�w�<�I�v�j�QPG��(A2�G�R��L/^��~{`B�)%;,�N�������)�jV޲��ۂ%J��{���+D�5�1�N�TW�J��V��]T��1oe���^����DV�E�J�p4qFT�iW3Q��u�	z�&�nbz&%v�c�zCނ�QQ4� �$�mR�6���ő��1�Ի[����vSyG�Iگ���|PC�O$�:�Ę�E�^F��k'�Q:�%M����"	DR%g�#�� �G .���������Ӿ�O�2�!A�%�>sI����_��R��x� M}6�����`G�S"��2���$6���ꃂl,d����^XG�+��G~��N��H)!�#J��.ɶM�L|��$�2Z���������pMc,�������Qx���kHv�9��*� Ů���7�җʸ���'R*����}oM��t�\2�k�'�g��Z7�%�=V~�B��w䮞�
{�+���������Y�{��s�w4�דJߞ4�B��b
V=U�P�'wŝײ&�,L��4��$`X+����u�8�\�cQZi
<4�v)����Ŋ���Q��-����K�73��8���Бd����Zw,���!�C%F��V��Hq��2M�����@`
>'j�-���!�E:��@8n�Z�Z�3��0��>N�)A��Bej̏�N����@�Y���7L��Q�M�n����J:��i��}-���f%,�(W��THf+�C�{�m뢆
��$pk�����I}����ҧ���_�l�vufi�| ��db������ϰ���B��Ĭ4C�3���&1˥�A��=4�iR�a��Ne�s�:L ��½ ���[.�OboWg)��N�����%(6�����R�,�����*�}t0�^]�ʣ�D]t�,����ޓ�%�D'���)��yS����v��w�1��d�DD��N[G�+�͌�?���r��x1�/S��o��e!C>�a���JKI��aא�ƴ����\}�v����?O���ɷiaԑ��`bD�d��|��_�S�Rz	����P�/%v�b�z}w[t��3!���D��Yᰃ�f�{ym��x�:=8��@S(O�v�6$�Y!�$~l�FP���cg��ro@�Tj!�n��=��]|u��u�A�ui=��w;Y]�8}��6s������ON��4>��ʠ!��ft\�MN�Y���!����C��r@�1��s�i�P���4����^K�h$��1����n��m�XB����P#!�_7��g��ݦ���D�ĆG+N:���.�O��ǥ�B�)f��W�Ձ��Sҭ�?���`MZ���!��H��7��k�"���k��=��r�JX/�T����T�b���o[V
fj���k9VN�e%x�0�2G����Q'�^�踚�%�MQ�W8jT��(p�O������K�jƟ��?�K�J��W�/cT���c)P�G�Hd�	Wiv�X��X�NaI��{�PK0f�:�k	��m�u���l��l��Ş�;?�x?f#�r�;Ezˌ�)�L=��h�?w�-��B3�'y� ��a��T���Rz����UL��6x���^{+m��+P6��IR�sHlM�*麩�p>4;���^���r�^���܏&�3�>8d��k?&�����!�/Ǹ��S\-Ltl�bx)D��b��2�t}�_|�3����R��$�x(gBn)ˊ� ����x[�U�m�P�f81g��3�v;�5����|S�a����T�q!��p�l��Y^�b��E��C�I�poA�9 ���|:������{s��\ Wy˘rP��w� )��{)eR�$�E�/��	�)d�¾�����߽6[�|�F/]�6'��� yE�_ϖ���c|�^~D���5�L0�r�n������IT�>��P�/�r���ϩ�K]?��j2V�����iE��-���.6��Ї�*������~E%j=���*��_�g��f{�f���.5o-�g��h��<���
��9?hpH��ېL�����O��j����柯������y��gJ�%}@���NR���1�Ĵ0K����5���l&K��uBޏ�#:�ly#̅���<Qo�HrI�l�盦��T~\1��
��h�Jh3?���#�Ѥ������Ӫ߿�L+��ԃ�y����4^�_s|�q��Lo�a��N:v�� �Zi��b@]�'NL�TS�ng�.ͥo'Y���Z)�j'��~DL�Q9`İYr$�)�V2�fQ�^S��b��߬����q��Ȝ��s�/9���))P��X-���f���6ȕ�J�4����ǩ��5E6�:���62N'���Z���׫����}���a\|-7����:õ�����-�+"�h�>�{J�r��ݫ�AEnA�웷@��b�C%�!z��@=���(d���c���6�\�~��+���E��2����x������W<~�p6{�_b�*��y��R�(�dh���ŽO%�������ʅ���㨤��Mv�q�80�yH�2�����������3c\qi�J-|����3���O:���!F�������嬎�P������5�Oߺ�c��=?-�2�!�;Ś�&�WM?Iu�s)�g�=�3`-dh��ks@\�-�D���I����/��&Y �= ���"��3ۣG�+��P��������7���Y�>��h�������(�D��U�Am��
�A�Ľ [�Y�p�����%W�������t-����U?�����;�O��oO��&@�������"�6@�z��~�>4�����O���{ �9�ϕ�b��_���6�:����"t5���4T�09?fK�e�r[C�zA�,{����a�C7����Yl'Sȯ5�`��Nw���"�$�t��T+�/��Ր�F�/�grP:^o^��&&REzA��J|��&%��a�ݍ˜hb��ݖ֙>L��g^f�g�=��M{*8�)ΰ��x�B��W_���([��@hf0UO"�g�x_�6�uA�u�4{~��@��.)�8��)e��n0��ӂ��B���B���\��-��b����@��k�|NO+� #O��}U��?L����~�0�+n��������� �jS�U�A��i*n�M0�J����N2P�?�3	n����p�zܓ�l��7�L��f2�� O ^�w{��a�|-�
WQ�˜W༈���*�DOR�#��w��?�%|��^$�F�q�x8g&C	Cw�S�/}����������B<�����0�������~
��G_}�H��"��K�gg�7�F�	�]F8����c�j� L�Ki�ʍ.�?��jI�FW�O���Tc�E���?1Y��3�%�}���ɇ_�r]�/Xy�]�������I!�����ײ�~�^����`|����=��.̆�w׹���Xr�I៾h�= ���ݞ��4�hY�s���@��*e[e���WT<-uL��&�_D�+�w.!�zNG�(�d��J4x3��,C)G2�e�>~��E㫕Czܚ��ߙ׻������Ѱ�&�����ζ$q�7F��M���^�����z��Z������'�]��R�gYj�e����*�ߠ3��*E����������y��5���ɂ���U���\�%ڃ�[�����}��g+wG ,��5��p���\��S[�S�H�҈=~���2�ί�,����o�7�Ϝof]�)Ϝ�JE�-��By�=]X����<��"r��nB��4��\���z鼐c�ȅ��=��񝣪^TJsRZ��X�c�n֟�k<���	���j"�E�S׿��Y�g9��(�FX�?��������1�F�!�]M(���:�9y���W�'/���B�_MS���u]R�Z�j���u��(&���Ud�͐����������<4l������p%"Ո�r�zoeW�!�_��+����:�G"����_��ޗ�.�. 7��ً���!'jlJ�RA�Zk�d�� �u`ˑ�k��4{���Z�SFC��-��-�nSN+ s�I�Ɯ��O�w,�]~ ����a��˻��˝J�fnR�	�`+Q���'�GKR[f�<���흃^�R��0��~x���G���f���./��ov׻�*�=��a�]	�d4��
v{��	�fp�-�VB�-�K+iu��V�{d~8�NL>�m�-�/
z��������z׈1��6�@��I�隗�N� nH�+b�K�K�O�@3x�L0>^L]����������89��w�K$ө7���q6���꠾U�_W�0�9޴h|��ej�`k��!R���#�#+ų#�����W�P*T
-đ���Wp̱��
A���[:���ܯ�����{������&���g���E���
�,�a���oN�i��@J��aj��������;� b�Gg�J�^�ٓ��q��*j-��h/����P��8�A�'=�5�J �R�Sڴq1���{�������^�]i��QLNWn�y��#��&xd�õ-l�W�y�gY��JG��g@���1����><HָF
��ƚh�%��h���^F-n|����5�����XFe�m:~�[�^\Fz��+��%b�4p8�@��jG�����*�ޔ�����D��c��~(��yV�@ 2�}t\|�O����G������C0�c��8;3�3�>�_L����/�[ÿ������5�G�q.�n�!�5��ôg�YڪV���xung�u��R>�u\���8���B\9���V�p�/*��:��o�4�s�4�w�r��;,'���g��zD�-�9"����J���ư�N
����m�OW��n���	����V���=n����o79~���-��5����r��Q/%�������>������%�	L�����)��L����/������zfq(̮�l�x��n��(�N(n\��XYd�M�D��i���$���ꯜ�u~�k���gy�d1��*8 �p��	@�d�Hv�r-�n�q��$�.%���<�"T|�5kO����I_��~�������r>۾�$$}Q#����)"*W��s-O�oz�s�V̅._�dz��qS�~!|dt��8��w9��r�=�|��o4��H��ݒ-�j>-ܮ<,��;�#�2�\�Y���4�љO,��9�臭�x��������;X��}//���A�5~�'T0�2�"./�#o����ڙ���Ć�.A\�;z/F��H~,*�=.��}e?�������ۗ됷ZB݉er�c9SEBTox'�vϬ /�����T����R_�x�ŉrY��o�G'�u����6�u��_G�ncPV�ndJ�x�����{���:"�^X��2���1k���5�(^�DDNX@0�&�B�?��{��2�F`� Lq�b��\�L�Km;�"P�9S�4P��0Iǋ���)�H��,��d5<)�Ab��$fZ<���!�Y�e��t�^Q���Q4�vI��&�\��`U��K;����JQ��cnG?mo����M���VW��\bK�v����'K=����nl,�m(����c|�
�i��"�}�7����|`}h.3�u���W�WE��ҕ�>�8gs�b
�}���U�/^�� �>�l�Iuxk�PNÖMYxx��E>z�����*���[мJm����=3��,����yt���P������+9�\=XY�l,�{Ä�Ď�'��3[�bl,e�٬�H#o>��ں���͖=���]B!ζ�tηZB��������Z��$�07־������-R�}��·��`l]�	��' n�SJ��B�?�����	��U��i��s�i0ܗfF.������'��D��V����6�}����e��}���{S�O�9�,�����( �xn��_c�`��`X�+�3��5�TT;1E����sߤ�.v<#h�||�߾�<�y�t��<8�z����w��c8L�h;�%�GH�Hŧ�d�q�H޿�F�]�w�ź�S��G��?���Y.S*�.�(Y�v��}*W_�8�PkZk�I)ϋ nE^���N�w���_ǾŅ��N�"�W[�pYL��/�E�j��Geg2��nŨ�ՒrÂ��\/>�Z7����J�I��z�(�\�H�q؇S��5u�,Q�(���4Dm��'	��-f(� V��t���7G�"�����Va��0z]Q3�:�>�"��X��-i�:�(����Z�3i_���F
�ط����Ӄ�����էccq�Ưd=*�?X��Qx��=���W�3�����D;-�$��f� �Cb4�C���ϋ��xX�q��S��?Q4Ȇ�WT���~���������ՖQj�#.��>��'I�����ym�v��+Kt�	?�YΣ���e����v%�G]��t��9X�|yq�Kt�S�_�����v!��%�u�������ڼ���f0G锢��<�z�"��������H���x�&ns[�77��}*¾�=u^����|Y�Ċz`���R ��|O7�NVd�9���9�`�;�]}"�~�O�d�����7<��X$I�{Ra*���s�V�`�ڸ��!Ԅ�Y���~��7;�W�4J%B�#��4�`�����LS��p�0�G Г��4k�}D�_^�ʺ�~&�B(&L�>��C��!�V�}	>[��<�W�b���S�%s-��A��?u_5v2�-�A�WX��`�8��NQ��g�<S�ػc�[B��t��yxt�/)�k����0�S{$w�8�k׵���:ڮ�cJ�GĦbN�ϊ�x�x)���|]�#���$C�b�����bDk�Iuu�%%��	��>u��09�<��<�^gtp��X�-�7��$<��{u�֫Qsat�'��/�������K���oup(��?���p�$�f���kZ�;�+Vc�ۗ�f��31Wa�%��;/�k�2Z�,Y&����r�w=�+p���{�
�^~�6��B0����w��q�~�&M���J���HB���Η���Y&�J[(X�W�A�T��ŝ��8�T����*�ܐە��б�d��r��p�M����Tl���*�GvЕ�͎A����V�I=./#:U�j9��HnfJ��C�2�пa%��L�u�"�
%p���>X$%B!q.�>�O�\Ƣ,�^LSJ�X�	����8Top?Y�E��v�ùP�O�F�z�c��>�L��%���ӊ����	"���?Ұn�#���GY��=��/��]}�x�\�l �Ra�ۆ��9�����>�P1}e@P�6�4�;	L�m�F,sxh���i�R�L��^,��g2�s��m��j�zi�U,�����瑽����X�p��aÚ���R���6M7)�%�V4"���B�ĥ;�2$8Jr���gI/�Ρ�cKb�<�h�hfi@�Z�����]��m
�y���Rc�6���H�PK(��V����c�7���>��N���dp�L1u�&�f�)Ip[{�e�)`�6���(7�l¸��ح����:�����x�X�u������)�Q��46��/��H��Z	�����I��ݮ��஫(��������=��c�!���i_����j7D$����p 6�js����JsY�	��4�F�/�1? bt����D�9�eg@��꽭\��|	F8��2y�syp=�{��P]�곐��m�D���Ȅ��g{�/�K�cX��D��c��ITx~��UA��8Z�,�r��@��u1��#��W޳X-���a��UA�x\�!����'q__�������v�����g�����h-������T����hnOU������-F�^^�Q�+FY�ZT�	I�� ݸƃ!HS���������~�ƺ���J,vyw�����/���0Q"x�0���7->"�X߱��g�q��s��,h�(�cɛ���8�|ܐ�^�#H �*��~L��ӟMg;��'m���}Q���u9U�����I�-�	�ܒ�n�g��|{�-�*2�����%�2�B��(�~9|��뼓f�u�K}�O<V��i'>[
:E�^�R�^w�E��j� g�A�w{NH|�<�j�@+w��N���E�_Q�d����~~��5�K3�Q��q�]�L���%] +���w���}?4�|�ke��N}�]3W/�C 23'��C�/_��y�)�z�m�����Eݼ9��Q������E�막c�<4޵�p�X$����6�kQo�{7��d��) ��6�-@(�-��h�h	 ��+�������WU�Ƚ��k�C�h*䰧k�a4���r3�6E��[<�lq�e[V�:���$�vR-Ej'��bL��j�_-[{	��nƀ�KR�a��7���q�{X���xV��t�fֻmA�7�Q����Z��ʿ�z?uԙ� edq�"�('���U7�&��L}.E!��W����;�Ell,>�Ӵ��{o�S�UE����X�F��(�#�`dU;��יhT��ܱ�A'D��|O���T�O�NY�5[��2MQ^���n�g[c�~'��M��ݳ:������;Ee�_���7g��xS����u��=��q���ޅ\� �f���`:�&��Lǭ�8���C4��$ ���SM��i+<J?o' W�*{"K,�ZY����9�q�4��p�⒢9H�b���L��_Uͧ��9>gc╬ �hfLtgJm��jm���e�H]�P0\M�i��;j:G�pz1%�w��D��$�.��wU\�[����Uy��W�D��ݩ޵�6�ފ��C'�E���ٹU��䘃�������{����ʾ,~���9.�0Y�G[k���[|-�5܅��9.x��e���&��+$*z��
�"
���� ��#RM;����qgz�>�R�u�.�u�)��u�i/��iHBC�uDBٙ��[W>D�a�UrPo�_;�I�@|�� ū��z)�C�1���E�Se;�����S��9����a��{v&"�~��M#@0���coU�"8�����3~x��ҷ��Q�� rpb���zX�(H�I�f�����2�v�6\��0���;�X$��"C��DF���}@���_@OpD ֿS�97��F+��1gj���e�8��!�
\����`���A�~I�2�p���BH�R�)�O�/9��-��h�(P�	��/p�[~���{�@�,��yn����ݒjܧ�����['y���f6.��Xkű��En_���zY�
M�$��`S��x�1�C�<�7�la'��K<���[�V����v�|uxҤ���:~��� ��XcE�⇒�\��+JS�p���G1##�'����s� 	��eQ�,�L?�ۢ���~�Mh��>���U�8�V�{\�=/0%Yt_w��\Mh��-��⷗HB���,���[��pH��"!�)�-�`.�ho�U� �U�Q����@����ț�ZJ����!s�ly�	������U��I�%T8�yh�\V7�-^�c��r�d/���;Xc�n��G��?Ӎ�ĕ����^�5VO�����ONll�b�|��o�鬥Z2�����T��O���u�Z��	�(�5�U����srܑp{(�N�4 �[i���z��"�Y�Zht�*6_t>�?�Bx��39PPή+�ҰsG��^$5s2	�OA=�L�G'���V��)L�m��v���WD�V���i�e`R0�g���4�u��{��)E����h��|��}/)ĺ��!�D8vnAG���%0��p�B�dNѧ�f&^����BAץ�i��d���(00�9�R}���s�[sfk�N�_U&��������k]����:�9}�7�푇��0����x/���:ES��.x���"�.w(�Ҵ���:���3�`{�Vo�`Ovvf�S$�]SY��}��@���&I���:��yl����Μ�*ܺ��C#�.��;�օ��׺Fv��ƴ)�.����ꐵI����run�Wf�|յs����^YD�S-aA����͠��;>"�;� �,�J��z~h����v��V�Mi�pv��w�5���ǎ��5�Ef.��\�q�����]����V^m������W1q�V�ɢ�o��lYi��Z��[���,yR�1�HFʕ��,���.l��s�Iƽ���J��ر�����\��o�?��i-�I�����1=�~�P>��o]((A�2Z�f��yN�����Dw��8+d�;}�vV �B㽢L�N%4#n��U_�V`�����x����Խh;�|Q�v�&�W_���Πܴ�m�R�$ã�%����c{��#.q9//k����{in�apRpO�.���GV��;��k�G\-���k~[ZQ�Am�U����RUK�$����e�D���R�_�ֵ�M<��a�Hj�`x� 4&��LFU�]x裁��������y�.��î��nM�>�}���蠷ZDQ;��~jc�Z����0�:��ga
�J]��ۛ@kx�gZ�aϵ�<���*�Ű�*q�|�~[���`t�wxX��"Ks�U9�=/�^;n2���>�`�F%0����-�tz�B;�/���7���M�6��]�v�=Z`����3?'?�-�"���K����L�U�֟A����xj0�zԵ�?�����`�O�VVcP�-�N .a�yO0�
��"�4���0�J_��&� �]��cH�֨�{3����o'����� ���-����fPK.�PN/>�G�o3H�N���3�={[W7c��oqE�QF��o�DW7=c{��@vd�Ez�!6�_2��o^ێ�p�g�8J�_ȕ���,��
G݌�ŕ2/�5�����i7�|��|���}���=x��>�D���Y��DN��v�I�K8?�r�緶�½0��^�0�؏n�N���Qmz�t�n"ea��|��6��޲��7�o�R�.Յ�{����$���s�0�����˧�U�(9��4�rM�x�(O��G�"�5�%}��E�yJ/����X���e�����e���?�h ��ܱ�j�O���E��`�\�t�Y��|����1���`����ѥ=_��q1�pa�!�~����T1�U�dN}�e���G�G�]7x	��U�I�������cemna}ɴ��r?�Z;GM����71��6A�T�9��X���� �\(!
�;��j�Jġ�c���}s(��B;�|i���}F$k?��{�ňC�vԹo�1��|�h�	�Q&n,����?ȫ(M���Q�\�F�.���[��Gh�'<��s��h�\�� �>B��gf*������^p�&ט�&yN��Ыָ�M�\$� B�؛Ёv6�L��`�[��EjH��\��Ӳ��!bWc������W�H�G\�h�y��f���d�͑��!�yh@4IM�{�mH/��0�k��)��J����rԷ��6��g�J�&n`P��r�x��;/Iy���ԯ��'�t��5�ZԪ��$S�{�H��\���f�\Wk!�k>�Q�/t'Þ���U�{�Y��˫-��b`�}��n�]��}O�<z��b�*$�v%\�����������V��wi� ��kr2�:P��{�L����'����t���r��D{�2g��X�9k�Z��n��3S�3���"��U'�p�SJxfg2�� ��/��
��{綂��L�q���d܆���MfIF&6��F�>��W�c��
���!�'6����8fr��:,*��*�wdغ�C"�>��*3���sܱY��	���g٭P��r`^�o�R���/��C��;3��:t)�^�O�.n@������!U|��*��-��r��N�w
5��7c�j!A#2�y�2��}�@�L�-F�i+-�v"�+�m�#/NP��(j�э�<��X|^>�~���.��0�}�y����\"�mS�ؙ��eϡ�-�{�
���{� ��$ZкR�.A��r]ٱ(%m9B�U@;F��m)�ҩ�[C����QnT�i��[܍�u��t���ࠔ��יvO�Q�dK�����X�m3q����ܭ���M:���6��ə���L2���7��z(B@ݦ�%�Wd�֫��Ӎ���)p�����]2P.�S2b�L價y���������5�X��y�J#�5�1�0�>�8&%���V�:��P��,�qP� >�m�В���H��%t	,�Zw�^ \ l�w�~PEO�M9��*�H������G�0�*g�� l������Ls߹�%��[�O�f3��`�����`�Ba�R�0;���\� ܿL�g>��fU��{�Y���8��0i|���I��o8��*���g��>���oǀ=/-N��&�c��j��} ��)���^C.��@^obm��{�s��&��+$��0���4�WY,!R�ؙf�"��}��������Fn���]�_�]%\D�v4ߎ��O݆��p�^�txѴ����G]��E�$�L���qEc�;��W�p����j%�d5��jfu�Jw~2���΢�ս1��)��?wZ���/�q择� ��k�;@��a�Z8�3��8Y;l���4��ǵ���o�f�+�k��ހA6�n�F��w�����@���J�j��j�X��W��VdV��@P%��,ꮉi��VLf^	P�|9f��s÷��G�R�pƵLz_��#�+���4��yG欐g{�nsDOSi���G��g�S�&uD�U���X�Oo��&"WM���)6rV-&�#�9�ż�@䁠X䯆:tRZ-����q�t]�U��2�8����Bx������X;/Gk�����%մA�U��oD�C��g����
~�2���	��=�L����S�����Á��?_E����֍Qb��(O�%U�G�|P���7����q-����t��䜇�q1���?\�O�I�P ����q�r� �ϊo�Z���\�8��:-D��'mL@u���E+5�ޘ��fH�#L%�|����B��^A��jR��%�J�*\����r�:d�H�F۶��P�V☞�I!{7龡�N�Ti�����ѝ:/�>���)�KèT#���Hk^�,��S�xU�&zrL�G�|p���)��}��}e&��43���SX��s��~"�'����rI�>)X��6G�̇0�E�����k��FG���^|��.Vvr�R�A��g���0��Rϋ��{����;��>�>�
��L�xTW��V����goQ28R�� ���1��	/r6����U�|A�7k׋gB�ܒ��$y:�=^�D�mm;��_��{|#Ț�Z5�m�c5S,���>/�a]�?Xb�E��b�x��_1�\���Q��4"��޺���s�`D��<��E^-*yDYӵ��U��0�q��`�j[[<[G]<]}^��gN@JH��G�p��Q��قX�����:7T >p��"��)8mA��B�6�0���^hKZvB�&f��0,�:����u��L�|�WѦ��6��>�el�iG����k�#�c��T�S<�f���y1
p�d�� ۱^A�R#�vnq3�Y�.C ������_^x�������%l}�(��n��a{y���ǝ00�^Y�W��Grk���ҷ��>P�٩�yi���3��u��.fPn9���e���D�G�ح�vU������^�ڹo��� ��i&��Gߔ��==(�C����aj,��� q@���0A��0L��;�(?U�����|gTd���b�������)N��AF�8�+ǐH%����zs��Y�q�'ì/�8°�]Ĳ��a�\��J��$��xC�Q�KX>�Sa8�Xb�O*��ۃ�@z��Y�+��QE~�#�s�qD+�@x�B�%G�S�0��4�M��/��
<y�i&�����ax&�`8��	�r��?�>�_|��ϼ�&�p�	ބ�� +���/!�]ӉB0,Н�\?�0�� �L!�M�aa�D6��͛`h�w�kTNak�*D�����"UF��@W<���A���JF�i[G�\������X_��k�=��=r^}#*�)�V����u�T����[���o~�+<{�>������%!��/_�W_���{�����轷q����W���/�P�W�B�@������6���J��w;r����ϒ��)��t��S�$&ĻZ��Ѽv>+K�V��υ�c/�;.�����:�`8�0��s��aI�&9������
�`8�0�UK�,�k�e��Nk �e���q�c%f���A��ŋ|BF�%6�J��h	���Y��X°��a	���7�c'�Jr4"-��ҡ�5y}�.����S1��޵�ڀ��E�;j`�m�����kfc�EI�T���Tw�W�Wy+"3�Hԗ��j������ ��a;�o�;x��kÑ���rt4:z122���~�K�w�y�t�5(�e���6y������oKA�ހ��^L�Y���2D&Ţ{�O��4���j	�Z[1�+Ga�#!�R�}.@,b�T�@�x�ev7g#;@�۬�&�s(��$l�@�Au�a" �@q�U[$@���/ �E3<�E�& ϔ��^D."wC�)W��������1���Tt���3�0�b;�t��x�n��.d�,��L�/Y�^~�Ë�����d������އaq��h+���ko�0لp��ks��#x���C�MH�����{�A:�e��j�ڭw�C(BDd"�/�{��]�.@b��f��΃�D�̓4������;�����%0\�`8�K�� �݁W�]݈%G�ې��3�B���;�A�Ώ4���FQ>�����U��s4�rEe�ȭ��픹��h}��	��ky�fv�m�q�፤Q��l?
ó��������	y�	��'<����?�3Rr�*�E�4e25y-:�Vྦྷ����7>�Ͼ����!�}��}�/�{�Q��C�����X"1Á,2p.�0��!I��X4��M�>4�l��0 C�K�́ޔO�,���g4 )ь�x"�c�$��Mu�������F��箆6�	S�vS���T�/.i"������:h󛀔�h2S����dp%)ըPj5IQ������8D�� ��KL �� �Clb",.';������M��L���_n�r��t�idf��f�!�����X{�8��0��"t,\���[�-=l�sP�܍ƞ���#,+��L!�L���+�]7��0<��I��5#,��l��iJ%L�pX�� ��A`x% <�4׿g9�1+�a�<WV5A�m;a8�z1�0,�*ff�B8�%R��$axՏ�0�Iv��{���p!���@pH&��aA���<��R�V����	�齃Ꮞ��@7��K�i�wXN(�辐�|v�� ���0�,axd���!�$��&������-b3%3Ν�F�Z6+65o�h��al[s'��\�u6�%���D�OFs/��x>�̢6�0�.��g��a�����V�~�)�ٵ(�o��Y���Z�'�=0�o��%y�)<��5��oÿ��G��۷��_�����s�����?� �{���Ky�5+�	�(Y��a�S}[���ݩ�库@���;��޵	���|��j��%?�Y�;v�wCG���v³�p堂�d�S��}[�{K��V<��Q"�>�C�b	���x��X	��P���7Y$�r�5���-������!�aL�FD�s2|l���9�'0,�x�M��v"=�����-�&���j��>��w�|����#��������it�ma�]���A�����5AÆ�J1�#2�ZK�n��x�/��O"�o�ţ�-Ǌ��B8s�p�����������H�{R��#�#ς.a.2�"�����e�i�!�`c�N 5�qH�J���i����x��c�!gX
�+c�t�"^�g` ����j$�8%ũ�aaX�n���r�SdP��JȠ��v��$>w�<��=�a�2q2�`��)�"�A��<�2��̌.!�����.dp�Yҍ��*�	���ݶ��2���Kp��f��f�߯��������6ӂ����/��'�����H�bg���c�|�=#7�FURZ:����`���'�c��{q�d� .%cKW(���	����<|��F����زe7>��K�\�QIpz�p�#O��COAk�#&E�-�]�G�<��df�e"E:m�c���h8��s[?��H����L�(��g.ꃣ���XK:�[?ky̥���x�#�Ө�X
o+;g��UȔ��2h����2{;'ka�Uy�C0�lQ0�߷�$�~���a�I7$�Z(L������Tm@V�v5m��q�A2
��41v_~�z�q<��s���gq��`����$p�A[=-���T�Ĉ�bU:-��i0W��0<���	$�GLn�X�򐚞���|hP�앬+>��Y���BzZ.��i8E���0����g�#f��1vd�����Ip#35c)��*�-%��LX���MOcr�4F'��D[O3�{���Ӂ��nt������T__�RWW��h�V��ԏ��2�4ԣ����@�0h�L6s/6pi�x��Z�1���".Ë$}>�4n�4:a)D����q��e�ic[Ҁ����j���t�4A�s���v �mH\��:7��Í~Ĳ�Ĺ(w-���S`xIe1�ތ��F�Y�c�a}���,��M�+_���=���C#&�|g,���taNv;���ϪD���mu2��U�!�bR���αʭ��R��K��QН���a3L�<�&I��f��>5�3��}�x�%f�8A�/ç�`XN�`�������	������/�mt|m�P2���Z�0�G��� ��mTR0�'��S0L�6�R��Z��zj���(6�̈́oS���!�u5����:��>$��+��h>t�C����$�E8��#�}9J{W"����z?�g�����x7�z/���N\y�-����p��7��K�T������#x������7�o��O���_������g�������_�#>��>������B���"�o9rzW�ݱZ�1{�B�(�j��f���r���lm|�֮0v��BF�Ne8[�����a7a��ɢr4zl��$�a��
��R��"]¯���S,�Bp \�Z�J�O�P ˺�_H�D@���̄i��[�����ya�{�l̝���,�k\��Y�C�	��7m�@����Z��D_4�$GL%�(hZ�ʎ�(i\���i8K��˕���%�6hE�4�Z&�׸��K`)���S?�Lo+2h���za��F<a|��Ƈ���/?������m�c�n\t�UX��\��|.V�ٌEc�(/����>=�t�2D����Z/Ǣ���X�Sk�`-ao���n�6l9�\���=x�����[����	YnT.�9�1E���#�X�$*^%�/F�=����Q�tgￅ`ߊ4w2��/�H��#=�#(�@e𙜐 ��0%��0L�*	���{&̈́�h�tSE��4.�1̼6ϟA���O4f��܃�:����"|�����/`���Ѡp)�~�#�as 61��8t�%�ܳ�&�
O�u��������62>&��g?W�Ϛ�lB�%W���^�>����h���/G][/"�a�)�Mwޏ�o���s"	����1>��av��G�⚛�F�ք8���]�ٗ߁3����.�Hi���5�݆xW�Jϔ��AXb��r)P#c��c�y��v�����Ĳߤf��*b�.�!O�ٴQ,�b � )���q�.�M ��6��y����Y�#��lR0f"��?hx���pa�����.���?H��#�R���I��E�0�g��D^�@n�`�����M�X4UcȬ^���F���7�3�AUëQ>�zv��l���(^A}�j����Y�`8��%�ASJ^#N�y�'�T4���a�����g�Q��Ɇ*���Q����ӘΠ����s*۔���J�I^�yHb;��/Ed"�S[����!?R���]��{/��)�~�-~��%B�8�ԋ8��Kx��cx♗��/�u��Wp���q�ȳx�����!�|����/��#<��_�+o��7�?�s/��B?2e�����+�b$��tE��*D����bDr{6���~�6?I� �T�֣	�a4�EH���ks�]�xG-b�h�m��1�jD٪0��#���!�aɄay?�-�48�0��9�0��z 3���C0YF���/A!x�w g��0�Ҍ(K�M�Ȫ�������|�勐(aT��,S%f��֣-����é5+i ��\�%��t ��N�a�cV LE�Á<Ä�a��^�5a���*u�x��?��/,q�6��cM��b�τ�ˉ�����|����կ���g_B��U�i!�A��&�K���.x{�aX���섶�u&�=�B�� S-▵3$���KL��Ǝ���}��렭]��҅�b���a�,�x����"���`���(�^{uF7��K|�Ͽ�g���x�����k��W��[o|�w�� ��_�7��_��g��������믹W]��_{)���2j�rl۾��v�zYw�1�� �Ok��M�t�zZ�z]�h��q��`,��`�|�K]�bh�H/���Ȣ����AxNc�uax9,U�0�Vg�^�M��&X�X��g��f}����"��z{�X�_Y�rh���N���g�l2C��AdX"�a����Ĝ��G*��N"V�%�8>'v�.3}�86ƒ!�5L �f�J3�#��:`(샹��Nn���|�!�F2	��6�!�ӂt!��GA��e����o���O���}�=>�6�|���x��Wx��O��s�a�eף�����D���9`ua��mx��s8��k��ѧp��Wp�]���>�k}D}�7�����>�4�;:�n��bHM����a(%$V�Cc�e(C�� ��:����tG_a8�l$�J؄����ߨ�Ql��:�N(�Pq�/�����4V�	�ۀXt:�$�K�$^[�i��
�s�!i���j�h�yW݌��z��M'ΎNAc��?pS�w��v ˒�.���Ʌp��8H�#���<�"�\z=��t���[�y?�Jj��y�h�a�%:��$����}�x���Q�Ѝ�	����@� 뗻�]}+n�� <U����ʭx����Y�]E���aL�]��k�a�་���o}B������D��k
°�I��Tz�xoW@4�d�Z"�wR^'�sB1�8��w�r���V��Le�;���/��q	沓�t6"�|>��!�{
�.�m@<7�M#�ю8v�1�zv�4��0�^<�f���,>�º%�$�� �pa8�`@�@��]F�&,#�
 ��3��I�0,�O�0� ���c�x��L�gT�XAp�>�h�����-B|�$`�2,���o|�4���#
�����!t%H�x|b!����4�Fv]�4�S�T�̭
�b��|�4���%������A�q���	�4��g(�Ѡ�ϵlSK{�Y��᪆��U��X��&��~��;/����H݀�{o��=�+m�s���Ͽ�ۇ��^�M�^�ͻ/ö�W`�W���Ǝ��c�%Wc��b�΋��1�=�ə�e]�%�Fg��+E���r���
�U0��Og����c���1v�^;�18��q���k���:&S���c�m�B���L</�M �����gk��$�W�"�f!p9���Tx�|��"0��{����Q�9����3��T#��H����a�@[2��pɅ#H(F��g��p���苐��f{>�̊�HoX��ڕ��pa8�4>�g�0G �#�b���`8�|	��O��þ '�S����a���*fX�$>��K����?��σ�����̈́a��p(n8�3C%���� �+<A�{��0\8�9�;	��t��`8�!�c °���Kܺv������aS�:��R��v߻֮M0��Fv�42	���4V��v�>��AO��"I�8�лj;�x�9�q��ز�b�Y�6�ƦM�q;��=J@~��K���q���l�R^O��h�&H.-��n���[Lظ}���x���{.�C;�Zvx�t��[F���"<�Hs\��r��l�E2��]}�q�!����Ԝ4��	�]��+g�p!�{�-=�,a}���,������x�ei5�����t��'�Ń���w�7���Pvr?un�[*$uOdD8"##��y	�8;ɂs4�l��UXDa8�"iŚ���}|&.�kN�
x��^O�B��F���
I=7�/�C��q���p�.��j�Z ����^9ia�aF;�0F����q�t�8��x�����{_qy�<y�F�Ӹ����qխ`�נ�}>���f{����J,X��\};���^������s��8���p�u7��[n�%7܄���{.���ٞ2y+�E�c����]��ջj�f.��]�$~�uTAc������C��Zo#��\j�dw=R�ҡ�DOB��'�2�ZH�"�
�j�{�g�pP<6��IΫ�D°�K/�&�s�t��0���i�8�
�g�������P�;�u��@y�0������U��]#ː�u1�rK[�����9<��D��v�W�#�:G1�R̨j�5�=��nD&���,!��ź��U�g����yJa��\��6cz�,Y���Jdي�K�z�E�!����[�U[.Ds/x�7�R��[p�e�"�Z�s�MH�;J�4Q����݄KH���&Ȍp�`�$�� �}|5T��`�+(�ߥSn�n�y��F�p�Y��7�bl'��iT.ڥ�7���loż�:a8�l���L��ǎ>��p,�����I��>���y�)A��-��&�2]@��0ub湐�3�0A��RP�I�ߵ����uT�����C���X��xx�*1%�W����In�
Q�o�8���C0�H I,YJ�@b���q��(�o���0�����T?r�(�7� �x@q,��,"I�'�e����\��簬i�F�4�c	��,�9-j@����Ɂ>C�Y��H�"�!���m�xo��j.��ꦡ�(Q��L2>�54vپr��">˃جD).C���XO`Ϯ$�Wܫ	��Y��{�d9�@�E�h�y{`����y%���Y��X��Ʊ�G�	��4�A�>�P�a����m�"h���G�e2
�԰����?�����=g#AB��$v�+a�Y����$'Iܷ��x��g���"����_-�J��X*��MB%b��a�l��U1���1�0^��r��`��o�53�4>�B`�#�����8$��`x&�I���K|��g
���/	��N�p��j��&�� �&���0��*�'<�
~�� ���m-LA6ul��{l23^�f��hY�5�ô�iS�BQ��������T^PKMZ��Tt�`�'H��IY�X�f�{�M|��<t��+���\��u��T���U5���GUZW�ڎN\�?����q�W�nuB�·!Ǐ�
�<��"������vBAE����u�@��A��K�� r
�'Rq�D�UK`��6u����ak��a8[�Ic���)��ez�O����w� ���E@Y�
�����9�WB+N�U#�<̒{X&�ȕ隹Oh���J٬�a�����aa��9��sRl��<�4�f��:p3�	��|6`\O%T�JU.�l���Oo�"��G�W8M�
�x�i�p�ܦIx� �q��8�Br*A"�����`م��|Bf*	�mQ�5��e�02��]c(��Ga]��4!����)�dc����؈��*�_ъB����6.[���W
K��*�1�ւ2�������) Nf��b,��D4��\�c/�8WM۝�(�5�i?��&P�F����l�<���y��&>K��������aJ&�(��ڕ����{����:y�4�SI�T֯?��Z�4����ۺY�����cM�p�6/Ca�0�2�f�A��q`
���63��𔶣�0m�������[�J�7oY�%Yճ��F� �&!�Y窐S�	#�m)V�3l���K�j*R�市�~����
�u���9���yj��,iELf����Uދh]!�h�$��M#@��e�@�&P�pe����NnWR
a8��?$� 0;�Sĺ�`y��1q,�s-5Hoq�Jx:W ��]�]�.aǶ$�܈K�_m�r���:1G_�G3���e�����q��ì{)����:��[�~�'����`�$��WtE��x�EI��E q�x�+'�R�!�'�����R�	�	7�!N�/��9E�s��&E���|֔,��~�!�x���p��F&����@B� �/@z�2(-a%�dҸO"�Q��0V�#�t�}%�M�A�8g������.�����P\��b�]�|�HBr��y4�J��2���a�J�ARF��Z��fiL4f5n�k<��.A���. ��*�����z�|�L�0�A�#S�'���П�{���b���{]T
��f����&��p6�C�%�+�S!-?�a����R0<+�Q�u1�5���Y����ʑ��}f˿�%c|V}wt�7��ᳲ��a�q��r�2!�㑬o����0,�#	�s�0�r�PN6#w-�E���mw�W1ÒM�/�R^�>��W�a��t�p�F���g����04�A2+�_���M�������B� ��2���3ZA��1>5���0�`X�Ö�Ͱu�	�n��q9�i�w8�0���Q��!��pA4�V�h+��Q���J郖J�:��ê�{��+ᕷ>��o~�/��>���x�7p��+x��K\��y�=u�~I������~��<��KH2ّ�̅��d.��ٹMT;;�.�s{��e�cc%��^��O?� ������	8:W󷮆�{5�-���XW����d�-�K�3¬'�fg!;#ZM2*a1�-�J������h-?�wX7���̈́�>�y�^7AW����)(v�uV5��l2�$aZ̋�Ysf��h�N�������d�ec+S_Z�	��*<B�/�r��mU�l�|V��6�	�^�V��]�m2�.���[̊�
����T�V��-�OP$�y��y�eCJ6���iQ�h��
$����.ⳮ����%h� �̜z���Y>*�/hB�'=a)���YcG�!��<$s�u�@�-�!�����4��$��b@�Ƅ��P�G��B��ʭ@y� V�Kן��+����Gş��Ko��_y�Oo⾕0���]0��QNk��{1��F���o`����"-��P�@�qz��p\�gK(N+�h�SK��bѿ�O�a�#��S�k���+�`�B^�JW@O����ae,��;[�L%|�|���Jd� �nH��$��4���y��4k�1`&�5-����Y>d��Q�6�W7L����|��ު8˺�1)�r����;#�����b=㻖u9p�m%����!FW�����wa�2n���g�(����h��2�v3���H`�L�ܽ,{ҩ&�X~�.�E�3L)��,�3e��	��رw`;j��X7����2Wa�Q<�Y7ɲ q��O	!�ނԂ~䲽�	f��oe�;�3��ú�ɗl�����	����U <S
vC���&���+J�6�^Q<�7���������v	�PL`��0����D��L��L�R	eie+�RKW�VP����R	۩��N�X<N�^�nK+_��
�K���˟��3Ʉe�yMSJH.%\/@�ϔ�Q��-&@#���,8����b
�#�`E@����alkB��Y����<�4N�`a9v��Ybx�r0'Ջ��B�p�
��W �0,��°ԧԼn���Q��ƪq��!�׍#�K
�X	���Y�e0���x�%�o8a8�0����" ���Q!&I��'`X�"�KWR����(eaf9�	��g�)�`,�E~�$�'m��O��%�t�'/B�� lj�lc���\i���-�k�>�|'����eD�MG�=
��a��`�$��"A8���L�	�!���1V9���$n�P\��z��:�ѷ�~���C�! >	�_��/>�Ͽ����J�/\��/�0�G�D ށ���1ç�$�@X Y@Y�²`w*+ ����0�N�J��0l��B �+�X�0x�y���q6����) NcHeG���-�]�w)2������_��[�PӹKV�G����/��=����
o�~�;���>����Wx�����=���x�_��wq����yPs
a���U�
kI�ŝ���S`Ƃai��
a+f^���^d9���бRgR��q��r����ѽ�)��V�I@L��#1˃���:�	��tғ�IID6aX&�p9,j�9AX��AVF*��Ttu��X�Vc&&؀�^�c6,zn��c�\��t���,F.-<�ٌ��LD��bNTΎ�Ü�d�pNz�J�l/�i%�D)��4O;;�>�@�J��E蠅N�M'PX��+��x{㭄%W3�K�Pҳ���(XBi&��x�D����y?J:V�����|�ϒ�+q�2�����R:@��Ba۔�1�W͇�b&~g,뇡��꡺pΑtm6������;m:��&6�~����a��)���b���Rʏƾ�x���x������Q=����>ƛ���[v�< NgU����w>�m�\O�o@t��ϧ���P�(�� <�_�4�2��#^cb�YS�ƹ� �2��) ���'aX�,l���.h���j����1�#��j�bCػ��G�%���X�[%R���a�Z�����cG�/Fn�"��Ƒ�mB��Lh~�b��>v�EH`''�OFN3"���߶����'�ę	ێZu�G@V��N�;��G��B��v�:g,;�̼V�5��exV�Zi���`lz�� I%S��,�ф8°�H𕥂a.CR@L ��G�b�	���		A`x�K&-����!��.�ۦ�!��!W�W۴.v���lO|]k���N8���Ѣ<��;wA�׍��c�	��U�p�rd���O�aJ`'���X�Ϡx��U�`BM���SS�����`8Ib���o|���.Y��P�����߭E�J�^���I�|��{����+嵃����T\�$b�ƩE���r��pK��� :��*E�P\��
�]8�(*RT4F-�FY<B��r g{Z�?	���Y�3�QϾ���c	_��Q����,Aa8L_���r��a����FW��Ɖ��끎�^W� Y���k%�z�$�]
B��0Sb�Ո"G�ExU0\/�(��P�IH[$0̶���^��8�N�Y�s���l��"�	��8��X��a���D��k����}+�d7bvvU��I$�M4�Ι+�0�2!0,��Dˋ�a�>3��3�pl�YH��1U��g��=f�p@�I5���f��3���b;���D���_
'���$���dğ~�o>���~/���V�P��ޕ(܈��aX<��v�p�f%+e#�:7�Ѻ��e0WOhƑ%�-�S����4´�hk	T���*���d�TR�	��8	Y����iLm�[.�	�_y7֟w��k�U�_��Ԋ=�`��K1�c�ל���S��H�d/rZ�#�u<�T�bv^K	^�ȩ_�\�װ�S(n�DQ� o�tÐ�K f�g�w�,Bn�4���pwM�y���\3�dgRM�HҘ���A���sYЦ%#C<ÆL5�S��V�����"�)�� N#k`�J�)KC�̀ݘ�٨M�.-�,���8bS6aZmj
25<F⨭f�-f5}lr<��1'1	��fDf�bNf���]W4�[����<t�1agφH�%�E}���t�Ar�P]a/�,�����u(��@+���;�@�F �0�Z�Q;+r&��<�l��x�*��-ϭ/�#@v��go�]c9�=+�L����*o.�)�]�YZA���,#TU��'T��ذ����!V�C��O .S��{�Lfx��t����_aj�6�m�Q:�m?|�9�j���y)�(�k��K����?��`�(��IY��J�Y���R�Y%�K{U��h|MH+`y'��u�E'aX)�'ǝI����$�`X��qlN���a�[ ]� �]5^�׽�=+�a�!B��Y�hG���v�:�l>w��R:F�/��
:#M��*��g���A�ӕ"�V�UN���6S�}[�g�c��װ�pY��EQ<����G��8������~��WfG�f��d]]Bâ���s�Ze�IJ�4�}	)��v�,_��xcX��B�,�?�=3`8���x��4޷���B<K�
�c�4~h@ǻ:�I@���"�߿�j ]2�K&JV��d ]��a��Y`8�0�.0\������1�i���>�?8N`�T��s[H�2�F��$B:��8���$���	��UA�	��k	��WF(.�z�B�jj�R)�|�	���C*/ E��V��.ń��1����'�/��(�`T)���\�e�j���(��l�cY/�=�	�V`xnfb��.��b�
����W��e��ߙ0e�f��	*�k�F���S�����~��TP*�A���0�H�m��*eoP��`�|�h(����(��&m�I����p���p����o�1ioT�$fX`�TJò���	�Y���x��Ѐp��
:����f)۩ռ1�0,y�g��9�AJ�A����	û/�7݌K�� :����c�O�a9X�}˓}v�}|y�=��7���o���kw"�iA ��@���UV����M0S�J@V�V���[Բ�ƕ���e���"��?GYX���zd�6"����b��m�Wu�R���MQt�����@&u�^����ȩ����}�-�m���?�E=�j��4����(Y����P4���߻}[�l���g�z���g�{ף�o*ۖ�[<&o'LC;Kɤ�"���'��1���	�����m�ٱ���#e���i@nN�����q�f3�n7�n3)�Vm��{\x]&��'�%/z+  ��IDATϹܞﱣ(��%>/��N�ح(�PV����b�T���܏��"�򐟛���|�Ó������p�4&s5:6���!PT(�M�7�P	�k�/\mf^7sֲ!X<F�����F�k^������2���Z�+�p!D�Ve��y(v�By����Z���T>Bh�"�C��e��d�l���z:°���ť���p�t;ю*����(a'�U	�����
sI!���,G��H�͞l.%�VRȰ��Ͳf�+D�ŁKn����K&qNl��8+6k�;W�u�&Dfd ����;w�ٷ���o�I~Y�|�N���	å�a�a8�[��VEfY��AB'��a�+�$�p���0|f>�?	���At�
�Mu,��È�Af�lo^�m��jB��8"�Ʉ n���4�!^�,����F�d��d�ߤ;�^�/�������@4;�l��aِc�fW��)�ό�pä3���ձ�,/k�\�\^Sʀ�#��\��rGc)�����˵T�Z�Mf|��E�C�u4�A���5-O�+[mmRK��d�e߿G�b14e�~��\�;�il��z�e�А+]��v�����쀣	��W���%��!P��d_o ��W@y���a8�gҙ���u:�V�?�2�����J	���RB�,	�jY&�	��زu<�z��:j-b*�P���	�QAE��`+N�t9g�?a�� S�QE���� ���[\0��S4�x�������l�@[��=c�:'�
�X/��I�n������\�s�J1K[ a]�\-����rI)�0�]8�6�@�~#Lҡ�|���&P�(��iEC�"�F�_�&��ك0,��	K̰��c}�e�sʤ4O�a�)a8��=�����>�/}+昚�`?��D�^˾����S?N(��T���؊�Y�7�!�Dx��1��2s-۩r֛2�	�`���<���K��) �W���3�pT��	.�X�&@��ƛN�a�
� �?{ҍ��%f�p �O��'�����;'0<�& ��}�Q4���;	���۽����{&�� �[� ����I>)� pP&ʨ@8�A�I<Ĕ����9d��u*�oN�zv(k�+ak���aR�+�5���8[�b8�&`o�u�N�ŝf��]+��V�۾L-�	��h-5cp6M�.��);_��v����x�W�� �?���y4*r�7Q[���#�wl��k�����ȭFI�|�*	,fA(��\V!����]+;�v�v"w`������!�����F�j;�*O�^��Z&�0l�ϗCH����M�����ӊ��U��Əz.��m���ذj+&ưl�B,]4�%#C�[�m��׍��r��a��5�^�}��<O�
��܄ƖF8}N�k���"͝�9�2�Vt�Vu4'��B�kSЛIH0Bͥ0�DY�&1�y͓*s�L�!��"ߧ�?1��3�C/P^a���;W�{	+]����U�!�k��6ϛB�5����Kc��*�i8���	E�<T�����0��s!R���u�WO�������
��� ��[+��$��Հ�LG.�����g^���zD��0+.˷��+o�	��ى�h�s���a<p�	�{�q\��nX����F���9����^�qn���aX�߬�I�ocGb	i �!VRϩe��^�8��P��0,����>���9$�ī�����{��!e'������C��m��K@�c�H𴫑�zv(�4j��,m)R�޽���#��6��=%��I<�lS��G�x�k��CM��׹�#[U�� �t�n�_-�R@8��1���S`X2���3Hj�zp���p���jBj.���Q�*ƐY4�`��}����^�av҄sH��#�
 1�E��\d%��J��s�Lb�;�X%wmϙ���5�"����~u΃�@��톖���`�jS0,��e��@�<��� �Ј"��� )�3l8�����U2�� ���[B�(���P��s�����<\E'�C
m�B!1Ô,cOSh`]H��X��3����MP�P�����rp�h�R)� |R+N(�Lr�`8>%���	�p�KU4��8Zi!�@TLQH#+��ZQ8�؂��1���OXmU�2��9�k2�]���:�̲Y�s����'(<�� ,0\NO`�
Q,��"o���lɺ+mI(cF�g�|���"�1�Z��c�r�J�a")��e}i��g�~f��G���G�� ����D�VͦG�-�Y�.���%�G�e�@<���tuR��>̼��f�ɐ�Zh��AW6[�
5;]j)��� �`x)"�I��׏���ç���G�&�j&+��OP�ԩ0���0!���Ӡ:�c���$�n�0�ؼ�\5�ƥ�.��OQ�9H���t��aX��	�$0,+L��7���o��7_��_��������($�eP��ǉva�%]�a��TZ�f~  , �t-Kw��"����.�%��Hw���w�ŝ�3��=��ܙ{ƍK��!��w�=~�����P����~�V�,7��_�bT�	|_(�S�0��Z�d�o�]�s>v�ˎ�%KP���l}���5$^n�
�L�nk�wZ�%@�gR�7�t�Pea�g���5�3�E�M�6��ه[��v�������`��銳�G%�߉��cV�e�9��H5E{�]Wrl�#�ٺ;����E�l��fѼ�Ӭ�<o�	>��y{�j�4Қplv��e���@����s>��t���i��@VR{+k`cCѵ��	��߀�<uk�y�{l7� �)��gm�<ݬ��U�}'a_��W���u�˫�F�����k��JJ�Xvg��=�q[7��csbLMC��JF��Y�8�e�v�nhE{�/��)���?$2��|怆T�V�K�#SP�Y�y��{)+����N��$�6܋Q�Y{{!�a�|~�����P�~߫��~�rdr��#0L,%P��6� �i�>/,�'m���m�������	V&�t�S��Ŗ��T c_����V��{�c��	4F���6��vE���E��<7���qy�^���g}�$��������?j}65ZV���E�����`�G��u����w�-w����.��?�S,���~1R�њ��s���4�<�O۱�|p�H��5��2��cMUY��O�Q�CɑV�ab�8��Εv�����T����b�&J��8 \�WO������&�?ߣ�+Y!�gmE�gP7˘����7U��p=�վI����NZ�?Ԇ���I뭟]JH_O��E̕��N�j��@�ʙ[ȏzH4�[jr���#c%���T����L�O$����F3n
�W!�9�b����<�qӱ] ,�� ��P�W؅4:���5&�EQ�ͤ}�7�2%ySsA��x������nH�&�_#pmX(�>�+5\?F����?c����C̫�:�T�͸���;��J>�|;�=������_�0<#�� ̋����8&��h�㻯�b�1��<Cş_�aR&�\�����`�0DH��=��]�f�'�L��%^$%{�;M��Mwa�a_Z�077=u/��blV]~̜��;[�hi�h��y G&�棽�cMM���]?��Rt�x�4���@����ά���FG"a��	��	�����(�[4��d$�����1͐5�7���U5�R��G�+A�ۏ�k�^� 3t��x$̀�3*St�^���V�cn��s�������D��w�V2�\!���a1��+�lc�8`0�Zё�Vg�]��2�	Lx�dZ����bI��W	���r.~��2�~Va�f�̆�B���:"E��M�fc�Y"��6�m��2&�������U�j��6I��9�~��^�Y��i�Ti3���L;�~w��V���_�f�?�G��'����~۫�J;�H��I�6������(9�X�{.����R��2��l�
���|(NMƳ_��"��Yh*�,�J�L�$ε�B3��)�B�/$�l�݌�w����z���﨑;�Ru[�
�U5��5�^�
��댔����q,�p�e*�������F�����6���I����&r?��nB#��]���~M�ښD�H���I�Y�B@�Oʓ��u��o���onҐ�|�\��9X��,����`H�}+e�WW~y+��`�;v���1i��[	)��C.���~ʲ��;�p^>���+L�p[Jh�@��yK|�D�@����]/�IZ̮�}y�d��^�Ye����g���4X9��-��� �T�"��hV9��|�C�b�E��Wv*��Ox�U�d��L�l3�����@�Լf��3���ھ�"Y���/""iŴ)�L?��[�OL&��A����^�a�^r3��TZ�������{���zp�ߋ�u�_@��C���������v�B=3���w#E��I+�B"=^�������/�u�,c_3�X~�v��#ə\�/cت)QZ���=3�0���E�	%�0k<��]P�q���3Ts��1<k�z������${���p��C�������["3\��浫�؊�{4`�Y~�����J��'q���T�5���E!���0�Np(�z�Ӫ{��jb_&'�N��΅3s��^��(��k̈́r�>�f�U�޳�K�d�t&��2)]\9�z�ێ~9�k2���̫�Ƴ����C�Uvf�k!���J;3K�����*��;��t���٥5��Z�y4���C;��P��fsO��F�^��Yn<tE�5��G+���P�!���v�4e�����
��s�po�<�y�w=��]b�^�Ȕ���ϵ�S���@��1p�|���|����n �������Nc���XgPd�2�C�N��I����� L�#6�f�
�f��q�v�������H�~��@�}��}yN�&��"E��E��$��Izq��M�)��t��W ����x��P��:M�:�G�ޡ�.�����fb"��e�螖�P)��"���oy6+���� _,ŷw��;:��_]��FU�Rǌ8�jq��y�F+��h@P՟�C^�4��P�gذ��(�_���(\eM�]<�'*�J��1(Wur\��E����a��0�W���B��I|0�]L�Jo������Qց45Uq�׬tT��y6~!�A5>��W#�@���A��(3>�h@]#	7Bx�����^�N�[�-��_j��k�����if�d�����`%*ha��.M�
]�Lŉ�N�D�\���Y},�8���
?p�A~��;��ɐ����'��iw�{p�cQӓ$Vlǹbx�l�Z�X-�n���c9�yt@�\.�;�m�}���	}Wޗ�����B��:N�����མ�:I�U�t�����M���_�l}YƗZ�Lm�ylqP�U]���M���#䦡�Ǻ���>����61"�X���{mwm!�g[�(���Fj�x �����|v�s3Ŏt�\�^���N�{�xȗP�	��evq���{b���'>��إ��~o� 8��H�'�U/�SYN�m�(9�=�Y���:v�w�d%�诳�����U�jI�'�K�-1�����['h�N}���s�Y��bm�֧.^����@�V>�ۖ�� �����E�Õ����=Q��'��Eˑ�K}���Qts���/�F�|��g���bv2z��х���%�D@�ɳ��S0K�:�U ���<8V��f%�'�yќ�<��|�j��y��S�2_w�nT�ܞ�3}��F'Zho!]�p !�e�����TWwm/&׹�Q�)�cά���b�u�K���Y}�~y���_��ζ���v���`�n3U�,z}�9MW�4�ļ)f��HU����dO�g��=>�w��<~�ށP�kvx�/?R�|`K�~��n��=���[��d�� q1�n����X���Ox`m~*�Ypiw-�8�ˌ�O�#������p� �"bL	,P�w)ں�����*�z�}!h:�;"�4`��lO����$����{��T�s�i2>�@��M������`&����g�l�Lݧ��T }��L|Ӂ�<?�||ntxq!#�XlD���D��
�2Ej�Yk-���r�ۧ	��E�x�!�l���h�Ӂ�����#jA`C��B0�E8>.�?�-q���C���Y�'pl�/;r]>4������<~�h�A��,;�wYq�����Ӫ�S�oۏ�������������p=5t���i��M9n~^���T�~��.{����1��!�v��*��X�!���6d1�DX�����Q�s�Q�?w�X�j�7,��EAޤ�8�K�2yl$a^�(l�+�W0������W�tY7��"������P�qd���n��l�2FP�P�͋����Ub4�	������r^.��?��@RMk4�C�0<��:1�f�2e��?3`�9=�z�J��������:�i����Gb�b��d�,H��σ0Ϲ��_���?��(�N����Ƶ��!��t�/z�I��*k�]�����խg�7��͇]D���|m���ZAI
�E�@9��szy�e�v�������l�k� 4�"��Df$�������ZƓA��w����1˃5�ՍmwL�Hu�F�uYM���7_� q�t��_�QS+c9�s5����̈́��%1$ZՎ��'U�f�i��}f8Ň'��D�j��gH�>�;Q)����n�Ta� ���29��4�R(U��so��=ÃB,̆Z���0�4�c����/hEWf��e�vyL����?@�L�2!��Sdc��_�#Ok2�c�y�ؼhy� �1���{X��>7eս�6I)閒��33��)!LR�gm�F>�����\Y>`�Jy�q_�&�8a8Iz����M��0P��VH�ZF���9���w{)��%!}j��,��eu)Z@�ȼ�E: ��L��!}Ψ"����C@a����� &�#��r�6/	5S�\���v����.}i��(2o"�FF���ňڰSk[Um��oh0Jӂ�1�0���1G��=�����Ar��3S�،"6�*<iy5��.Q��� �!u�~c�9�ǵ|�����@���B��+�l[�������G#�]:��_z��N���;mbO�!I�E���Y=L:&,�3��N��(��|G�������Zצg�m�����^9���!_+͙V�}H���n�UV5p�f �;�0��x( �� ,���`�P�,�\Mc��f�?�3�CM?)E�7�f��*Xs�Q<[hP�������ʤͩ�W����<�����<ˠ���Zif%��?���z�����6�Ĩѐ�S�$�c��A�M����QS�s~@��a�q|�,�a��lvpT�YO���G�*�/���\���]�=!B�8g��|}~*EuJ�a��hox�>B�@/����#`�c������h�����2�tF�Qmm��?!�[_��Q.�����x<�]:��ҡ �f<�*�
aĊ�V�O�JA|�a�$��E��u�3%��퍊.����1Lb)]�<;	-;wF�4��KV��}��r��%D+�P�����X�0\�c~i|��D(��"��c�ꮍ�+3Ӂ�� � C�L*�o�j�-�\>�6�l�|	���^��cXoE�2}j���HT�uv�	f�=�\�!ӫ]E{�w�M]Ӱ+��vSqhE��:@;�w�����IX�Y����Ϊi_��(��C|�fV�b�P��Ͻ��s򾴘ꙮS�S�^����,>cE�n�@��K��ݰ��W�����yʓ�թ�jv�RtVa ��R�	�B�#�j�0�ڽ�D"Q�kq�P�� H0�"���H\v�k�5�*�8<��i7�y�~xT�-�IK'�cdg�Fޝ�qq���|���}ђ{�T�8�� &�P����ot��-�=�:��T�#Kn��w�<��Q3��w�3�d`>��?^�Ƀ�q�"��P?	�ھۥ�|�]�:,E�ֽ�(#���8I6�0i�)��Z��Ԇ��W�_�Gׂ��-�Ϧ<˾�sF�8{������Ȩg����؟��׼�
�
�l��Kd�ZgQ5��I��Br�����$K�jq�a7.����{!�_�w<6V3MgZ+�~�[�^E\��1Ɵ�:�opMf�͂�x��M{^
�|MU�Y2����N�7ue��R5�SM�7�C��C���<HÄi�	��䧲t���F���
��	U"{�
�e�Do";��މ��t�6jղ��_��q%�P�?�Fg`S������: y��):N�
7̸"3��0��4����� �2�6X�r���7p5R��P�!	�м�LD�0+�a��4V��	=z9�U&����Ɠ�Qݝ���|z��L��1>��`���/F#�"`��,O��~��W_@����p��:�+N�C�{�_)�t8�H�9�9_�&���`�=��%P�&��=9�l"���)mqɾ��*\�J���Iať]�*\W}m�����U���0=�n��yТ�r$�{�l݈��PZH�bf"Qc4'8�*v��Lл
�w��?��`��ry���Ƽ&Jh��z�(�&���7E��z�'��H�M�a:tFoÈ��W�xx(}cnr�.j�E{"��ͫV��I>_ �(�n��zH�
����/f�ょ�S����=��Я��`�t�<A�V��`P��B�n1x��-������>��������r�x�elqv�mpx`�z�h��=������l�li�������ޡ}np�Ʊ1�� �@h�N*�Bl�o�oF�nXE;.E���Py0�y}(�<Aid�����C<�?�άx�U3��Õj�^����@,����5!п�M��tC0��6{���dxuaKy������>�����+���oR�M?��gt�?8�I+�vO4>�[�{?R��>�����'h)�f���җ�p,
��%��ݢ���"�mb���0�8`�o��b���@c2l>)0|�TJ1����_JypSWڲy���g��2e)��e�ۤX�5-�v����#U��+�A(�X�E0�T�7{�ȳ!�L�������6V��?Ī�-��K�$E�'�&ׯx���X����)nrS�!מd>�����֡B[�)���
q��He�u��fp�K�+
�˹Π��}Q���g���؜N#�RK��r�Ӗ�Lf�zժ��K�BX����ț��A <�����6}ఘdq�����ʜ8�����\x۞�)[oT�0��:�>���I�/�^�ɦ�a:ws�����]�xwZW���[y.X�f�k�&�ʚR�H�m!%�u���:�A"$��7sba�D�>�1nG���ì��ι�{������"@`c�ő�O�a�_w!yg��HE�/���x	�G���yŧ�M����j>�ԴN|*`@��������������64T.s�-�x�j��k�C��\n����a�6lB5t#�����e��a����/G1���ЮP����9�3��)`�0�.��H��Ë����˅.�{������1^�ON{Sr��u��Yev7N`3�3���3�^z�-bn�eg�����]�^YY��]q<(�w��7}D��#��j���ʝ�O�V��w~��so�m?�r�jQ��p�(��_!�g�E�:E�lX��ẃ�0y����)�"*�	����p4��G�Z�=�2ݞ�2f���G�-^�N똨|r6ZҽK�q��H4�適E=V63�0�3�́��ꍨc+ii�#�Iڼ�`�]@�� H�~XDO^=��W[ƾm�w8�'�<p��\��Xʝӗ����h�Z����c����W.�T���F�s���RH��qw�D:j6�A��5�D�� ��Q�3{fw�`i��60r�~�kYs����=��y��{A�ˮ��7snWA<��J�/�(g-�;����h<������F���4�;��IxCL�p��q�o�oޜ���v��e�@�*����˽�HA�2;'>���6�kf��SC��l�)�ۯ�����H{��cI�h��B����-�q�}k�d���i߆�����[z<����ō����$.��l���\����OJ�LXX��*�}�|10��1Dr0��b|�8��X�����P��r�K�1��`�+r�󒺈�r>�Ab"\�A,�iF�=�ƽo'���N�C��v�x�:��Qt���Oj�Ռ���1�OD�T�X�4�2?KZ����H|�I!\����}�&O*��܇��(�k��CTN�%{����فk=�uY��|��{]�|��&��ZU�5��X����7��%���U)�ٵ��L��Ӫ5��{�����֊x��@��-�=�:h8����g^���D�"2$��&Cg����t̟S��C�T
S����e�!��(�D~����������쎧��擐5��� -F�B���L'�������BH {�4�>�e2C �����P=r4B��1
��/�嫍l:e8Z`��V�>�<����0�>��j{��xv�{�:�8@�:}�N�,T\|RCژ�o��A�.bi �>n�rę����������2�*4W�ط�Ϟ1�I����n74�<��>類�$�;X9s�	<�`l�u�`�`�]���W~C<��6�Gt�����^�K
'����w�=��!F
KN|�s��k�&�t�<u����"��J�X	��`<,�>��X�*����E��[r���m�.�)'�67x�^Dӂ�J��[(e����c�>\�.WY��2�0��F��0u�o�!#~��iO�k`*�z�-���Cb �U��[c�!���E�U���}�:F��k���+�ݕ� �^�����	z��|���*������	�Ak��>�h�+J:��hz��%δ%�M[�N����e��*�a����ب23i�{�SkŒ����f��Vf���o���Ff�2����ּ\�*#\y����r�wY���E�N��~�Q�{��gk�U��O�L�	���Fn:>��L�\�?+��5@s�~��l^h-�!��r�v��h�I��>��aH�<�ICx�1�����%�v�zՍ^/x�-],3A	�-�;��H"�CF��=���������1�0`�u~Rxg� �<�s��b�#!�j{�)J�p�H�ٔ��㌪#�5�@���$�w��i��Jk]�v�R�X���&�O'�+
_�<k�|��i���m<�=�RQ�p汝\{.� ���+Ak`fgϤ��^zEz9�<�-7��8w���uGq��X�P{^Bv8��+�xP����������r΂����4~P�����n�L܄�x={8�9Ӗ��N(�՗��t$�ݡ�UD�y��o6"�t�!�����V��5���D�|wm�� ���"7���Jy����B��F�/�L(��v^�v��O�I����O�<�ظs��볥�%�s� �J��ئD/EHT�:hU`��V�>�T��4n�ev����0��-�ߍ��;CD����o��b<����z
��\�?��]�4|��f��c�.q���G먠���S|H���҅^� 3ݙ%������/��H�H��#l%Z�J'X^vd�{�^E9�ʣL��`��(3�����Ds�ط���5����8�����g.�(����q�󲀁��Ȝ^�e�a��\�o�S���OQF�^%��h{�G/���z���t��Џ$x	�zz����:Ħr�ʣ%T/Fy�7���u����	^�v���t`�Ƃ�V�Ox�>�Ԍ=S���?�A#R�1�r"�e���&��B��X��^�<SǺ�G��k��$��6ξ ��[*�h���"��4�MMR2���-<����O`
�盤��j�xGw%���B
�<���O;�#��_E�|ttiF:g�0�&��F5~��,�J�Tw@���)f�K�Z��4�A���%�. ��Y��O)�ʵ")Ҿ��?���M� ���,�W��� US֗�#_�D�q�IǤ�Q�ԞmF�m�M�"�?&���QLy��=�������/?C�P??ך�Bf�7�_w2SL�3$�Ԍ�Z�[��N��U
8̈́�MR��\L���Դ��V|�p(���]���B|����Ѡ��T�B��O�E��rU�����&�j���Z���}���{��w{@-�jl��ϟ]
�];���H"Q}�H�k�g�-ՀF�h5�5 �0���_��?��/Z��[�g�1���#��:`�Go�Um6�](�8>XJ}x�U���^�|�>�)��(v�5�HZn!�|��f���MV���&��	�K-^�/�ܹ��B��m�s4o�6Q�{))����y�1��Q����aE��+|�G�ot����������k?;~}ޚ��ĬB�
t$��fz?�CV�x$��-�{>V����EPf]s7�}l?��B	���U!�.�U1�4V��g9gwP�����|��C(�r�c`ܝ.l���W�D~>�����8�z6+�c��DR���f�g���f��7��b����
&O�厧�~�e���u�:�q(�ۼY�Z��q��΁�b�M����Ȫ�r�.���)�����8���7�*P�R��Yl{�à�%�ћM��*3������1�d|�����(�5���$��'��z$��r?O���w��#Q�F���C�h�Z�dS��$�1ƳI,���I!���Ss-;h��1����p�A��x	S�S��-[a\-G���պ	����+2�G���+J�3+�W�D����f����3��0�\`ۈ'�����_)�}�����͇�Uw�X���i��9�><�+?�!q������.L��tb��;;/���ܵP#��|��ⱼ���݁��Ǽ7��H?�}1;��q'^W�}� �҇���wI&i�.��}v�0^eW�hFm�eZ���,,�)nY�)��[Ԍ��HNEB�0bx��u����i���APq����q&(�dZAKIw�A��h՗����?�LB�ھ��Q�	bڿ-��hl_��,Ow��-��RD%6��^ %�E�j�[�fʑ�-ϕ��婡'�@��%��Q�/���I|w����L_�ſ̚�C]�e��51ctDR�8��f����f=t%3�^,;Ĕc�:����3���g�2C!�
�p]Z�1�=z�Ȉ���M�9M�H��X�:�����j=#�����'\=�y"��ف$���U	�x�pH�>2����k��k�jD=5����QFC�ÿS����HB1�B����!�o�o/�Έ3߳�����y!�0�A�3���Х"���P�e�ms2�t��6~�CrT������/�|�/����o��l�ta��+��j,,9��������Ҧ��_�B���SI�e��������%N�å�Si��~�ӳ�2���_� 8h)�]�mj�{*��d9��P��fr�s��MF��W������"֔3��)3%{�	aV�:���VI������O��%��+�S���g������c^�S��
Ml!�� �'~-Q���H@�o���Frd=�ēn=
 ��*
�=���P��Ϝ���P�@� �n9�����"Z`�1��ڥ.�Gn*#j �^�n�ı5=��#$z�@�,ׄsrBv�I�y��ې*���-U�/�E�3�ë�ps��|#-~V���#�|���kj�_��n���j͹��N��Un�K�0c�:�>�>��mv]�_���m)n�{���Z�l�{%h��Ė�|����Qq(�D u�^<j����������8��^Wg�?&��.o��5��V^���G�~�V]���rE�Qb�BlU`y��s�22JL�}�¢*>���V�	�O�k��\5x���a��X�<��Z��P�3��O���2I���̠�ԭ�N"bPP������Hx���]k��v�bO�1���ऺ���{���`0�Z�\)�Z!�@�1�z;��&y�1n/C����Ϙ��5c�S���w�{�}%Ǳ�0�ͪ�S��<p���آ>'yY��'�\�������?X���\qkEp�.M�/�8ꉃ@Lm�{R����X��.���c�03��4H,k���b���H'�k���J#$M�l$�C��s=(R��i���>W7)#���2�bk��TBqh�j�@]�9���s���K��gu4�(N�������*�d�q��fa�$�r_*��B������O#�r�½�r�\��%ӧ�Y\Mμ�(���<�9+�~�{sԹ������G͏��n.��l���l�:�-��]j�k ѶHf��~��`R���볐���IO<�F=�:<S�?�\mOH�n�;Rh?P�|�9�7�e�'��pS��g�iieg��[�2C8���� ����	��y0W�-�g�$��GQ�����Z�2��&
�Q�$/697�(M�B��U��ϋ&\�+PI���_��t9�oB@�����������!n��ƜyK�y�y��6�>�(�挡�/4�T�� ~J2&� �|�>A�8��A��:�\YLD9�l Ǥ��عhq�79%��a�P��$�v ����(�z���d��fLl���
��d�A��w�\[���� ���@l'
~_k@9�GØաM�l�*�^��8���Y��;>�?c�'.�Z������Sօ"��4b�XDb7��H���� b�*��/�*��@R�r-e�!D��es�'���`:9�i�~���b���ku�\��.4p5�5SzaO��qV�J��pn�?�)2�"w�E�T�!P�a@���a�ș�JS�É�N�Q|��n�ף�~=�P��%޿��lr,��d�����ĺ�~dc�.�8!ya?�9>���N�-@e���������g�9N�
�Y�]�5��E��l�����F�cS)�~ G'��6�%��FH�4��|pl���0��8\�@��\�=Ч})�_���L�ܳ%jR9m�T<���m�0���l���M(�Q��`��h����!M�� L�u���襍���� x�2��i�����u;���d;��o�pk- ��o���Ȱ��QbWN�#�uaM(��O��NYB����p�/�	�o�#�~@�7a&�NZ.a��#$%��AhL�G��U����'���[4���0SU�/�b��=?��V��	K�����*�fB.y�
�:P�5z�����-�Z/����8�D֞�'��A/���0�5�q�l��J�Y��m`l�@��N����hGɃ�OԺ�!���1�g��K:��s�wy�.�23��ըO��H���'�s�"_+�U�ޢ)�ɬv��B���@YB�@?;��?��V��/��b���,��i�?��j���@��I��V�0X��$��Y>T��')#,h�y�1ivr��u�1�D�$�vI1w)�C�
�?�n.ð�ceh�4 'Ȧ��|��X��`?ߟ$��1s#���ܾ�d��O�/w@����I���.Ee� OM����s&fH_>js�&*k1�R�����sH���r_�&n�=a}�3.k1�M���^h�┞�O���af�A�TR�#��w���I�O����H�q��6;�6�&�H������PE?�� ����4�[������c�������%�t����]dB��%�XxB�Rn?l?��W�V�7�Q�]��,G8�O��c�o�"�9 V�9`�tEf�n����X�e�D�[�EAw̿#բ�Wz��Z���/O��_��Y�R=Ib�]�>)�;�,�2��&�!����>Ԧ��w����W��!����1&�WƔ'�4�<q��P'�eh���"t�?\Z�N���j)7E�}0h����Ü�޼T�j]� }�����	�`j#k?p	��$�����s�rd'��j�Fzc�M�<�A)���Q]"&�w?�/\��sԕg:hQ��&��6�������? �֑-��U �`-��؊%�iٽ��Rą)
������렒Ֆ�긱��C�t1U؍� �����a��?d]�C��@ln��?�6aWQ���)=Zf+���V���b��;�<��`���𱟻���".�N;��q�:��Z����i[��A���	J5���O��Qk��F�XҖ³����\�jۥ��J��|�Ti�g�%7!�Iϊ��a$`xx�ݠJ��\.����h_)�����}��,V�4�ui
~��V_�ܻ�v��Acy�q���,������V�l[�ur�N�<͝���]�|���	��>�����}\^������3A�&a�1ET�s��_���9�����j��[�ڳu�韲�)���QٹC���E3���V��/��!(h��gꔘ����h,�_�(�x��D��f'D=}J
��	@J�3E��w��%}3�������ྪ�l��ek��k���0�����.�{�����7����v�����ң7�̆O��h��̕,��B��XJ�"�s̛�`Ǽ;�m@��ި���K�\�1MfLbx��J�
�X1��M��D� :�XEB�͏�
=�?i������f-�y�fE�u�%
"5�_��	!v6�Zȗy�{�Bz넲қv~ǔ��$f-��PM��|�v��G�L؎s!�Q�#Wv���
:���g�l�+ڹ�&��_�Y������X��j�p��l�X����2�m���Y�֪���'*y�%��w��Z��g�
Ĺ�<�D��Ǹ��a!�B�]L�2�6�EW�Z�����}L-2Z5�v۠��a����ՏJ%���.Y����.��ل��$�_�fK�Pؘ�Q���)�V�v��K���DO�+Dym��^w#BNIV�|��+�ln�л�m5��/�K��)��#֚f������(��?|����aN���� <��I��o�z@������~��s��0��Z�/V*/h��S?�W&�_�yR����+�H���i�u�w�c���_�w��/y.L�\��{~�]?G���t'u��w�*l5���W�"��1���C�H��w{�ԭO��@}���R�~~G'��0�1���+�+]O�$'���Ff�jJ�p����F�Ӟw�"��8HE#�`�?2MFt�魞���S����W��'��ڞ��p��?���Yp������L;���h�x�C�ƕ����>���S�{׌|l=�,���1K��6�b/o�n�W�W|qJ�4P{�ɉl�b�>��Vx�g�����v���ܛ�/&\�ԿgH46��}��I���8�X.�H!%���{�*�#��������⿤�_�]����3iK�sʵz��jΚ�Pp�J��|}�����ʺG��=e8��e��GTGp搟<�B҉��������E�~�q(Ez��X�zU4B�@�Rk���V|�?Nf�� X^�����{{h� ��t�º�i�"LC�m:U�GQ���A�ME���"∛�Hi������x7I�{��i#m���Dz�J�c ny� ӃJbg'��rΑ�cN�P���\a���T��c��(�1u�C�JI��xK,l��MF5�v�e��������S��3#�b�y�&���c�W��y��|!�hd	�f8���Z�vo?��B��<���'���Ņ�Reߟ8��s�s��!�Ҍ�S<AnB%.\��L��͟N��n�(a����Ko�AUIE}��|��YE��	E��m�l'�m���l��"���z.������*Ѹx�M��B%�5AB�z9��qli�9�u]4�����"ޖ�Oqa	x�?�7(?��L!w-P�n'��A�jaQ������;?+���U~k�_�
�xF�Eb��yŐ�J�F3`�rA��	?I^h�`l���/�̜��fF�B?�^5��oM�ґQ<���~D�G�^�9�@S��y�9�w�xg{���������ᥴ�z,W'�<J� {&����ΐ)�$��w_��34�`���w*�]���Nmo�`�om��0��5���j��T���S6�і��r��Տ4Q��T>����
�xj�hN����s�e����R�� y��k�˱���a��dB��y\���Buo����vCV�V�ģ���<1�Wm��y�_��u�	-�$t�֕,M�Ld����m�}���T)�T���N1}���j�Ė8�Ԟ\>�yO���C�ܖ�F���g.���ك�gD h�Q4��T����GA Ϗ��1IG�@C4���(a����,QY}��b��OH�֛=�+5�	-�/��Ge�/	1�(>��}����:��v������n�V�(fӾ��<��g��a��;O��/��}����$�׍�l��A���>�Y��-E����](������� {�[
p�e�՟�<t_�	��yj��S?wv�f��'��M�@�?b��4�o'���n�"�#�7�Υ��|���\�J'�؂���Be���Â�(W�T� �Ū�:#����z椤;��k�i�eU�b��?�y`��2|J��e�+˹"�M��S�?RX��,���Y��R�VH�c��M�%�g��� N@���yI͏"�e�`��*�-�FD�hD�"��KW�Ɖ�p��il��>�ml�d3.]8���7�����/�)B��y�`�3K���d�Ә�أxa�rl߾'�Ǚ'��¢��m����lG�����s�h��0a?�������%�}X��w�AA(X��&���v���!���
�Y����:BVTE/�ά0,�aI��-�e� ���"dhb6�b����E	�Z����Z��`؄���k��p%FL\���6�&���@s
�CbU��G@����	��&��T6��hj����:l�҈Q��蜄��S0b�T3��h׃��a��D�� G8z=���$ئf�����CQS׌���T���
���+�AnE���ZۀԊz��6�Z��UڌԂ:��r�g�!E6���*DHL˹�
��E�b�ǖ!�eHOO���G�V�]���\���[�waX���#�>�U���
�p��a=��SD�Z'��na�b��2���cAnM^ߴ��{N^�ǻO�֯��o����DX\6������´�������i/����]����V��d��VX�FASІ��gd�������q�v̘� #�'�i�pL�8�ä�f�T� 3�c�3<����:_g�<��XK0r�cP���Ύv�^���_|�9L�0�'O��o����o��3h횅�2�Ed�
߱�g?��.0���,?W�{o�Us9�0B.솆S���j��(�0�����0����m#��A7�ϼ��+�χ��o6�'~(|ے�ȟOBp���C:a�!a���p?���U�@8˪�L0|?P�V�?�~ix�F�'����F�?�j5�K�P �`�*�{�>Θ`տ#K>� B���O�ԭ;��3ߙC'�������#8����j�[�����m{�#���:���մ����޽��K��f��}
'/�����!1�IM�*�%�Ͻ�����zc�sRP^]�9����0m�T<��s�<q�	4�}�1� � �Y�H��Bay	R3�`	� %5�m�Hħ$#�l�#`�ؤd�kB�3u.���	�S�>M4�c�E�QD=#J���G#�A�l�i0���cD6�b���M���������~�
���{a�>�0�{�P<��:����P� �W°�0�5m���O?�U�����_$����;7�㏷��O�㋃G0n��U�@R�����O �VI�4=A�.[%aFn����j�^�OVy��E���W�q�#�q��;�Y���t�&� "&st�p-Q0������D�ŧ";�ŅU��i����^�PBM{�,Y�W/^õW��͍H+��=I�]���)i,b��^�AQK�|�^S��w!�e�$��<$y����\2	��0MT�6�O$�G�d� G�U�f�l�r.];�}��`��Mشq._��k׮b˖���xr�X�xV��
��O�}�O>�_���.�W�5�/^��{��tj�n���ڍ뗮���Ә:�	�I�f���,��0�/���g�QKH���Jh����&!0l$������q�j�)�~@g�K:0�.I&�a&Q;A�Ls�,��
	 K�&��G���?ˇ��34)��x}�v��	��=�Φ/�K��E�1�!Qp�7��+.^�p�	��o�|��5a:�<����u����[�u�|�ï8�6�]�hd]��=.�S�����"��Lp��o�щi�>�Q�?t'�^T��w��嫷�.R�3<���q����ǥÃ�n╷�����1	���Si\%�S�]*��r�%k	��	�/GPb%U�2D�6���
�R�~\��g�qBB*��X��0,�(*�D�p	ÒM��TСR�	���h���˭�b�s�TR��G��7���8vpQ��xN� >�w��#a�����O��7�b���HH��_�`��|�cn��~r���2����&�ڌe5�)��+-Ɔ���3=������ٙhւ�����>�EsGbXm�ڊ��Z���,�R���t6�`d}zF�aZg+�jK���)8���u�^z�9���c4;�Ç���#h휎����;%L�0^�N�����{a�D�<�� �p �7�\������:��Y��:x�7)y����RKUEX��gx��p�%"b���`*��V���K`�+��,a9�~���6"9����3��|Ц>j�>�0P�Vã��	0Lhß��0 �U�|H�"� q�'�k{���]p��PڶЋ�� �a��l�����๳���Bt�6Si � !���ɋ��`�m(�l���g�so�
)ipv�Øѓp��Y��{-�f@#���"*�
+�f�r�����(,���)]س�K�X�"�q�ڳO,~E�E�i��!܄��2��U�
�^���4�;İ��l�.��կ`<��;w��B'Lch�Gv�ȩ�8z�:�.~Y��y�%�:=C6��yl��`�	cfۦ�p��_B�1� �^��u��Y܃82KH�K>k����ðU6 �?�w�pBS��l�W&�����1ϭ\��K����[q�L!0|A�{`�? ��]a�۟������ѧ�`8q�,$���I�aN�����_��KI<�M�
��hH�`�L	�VYٶ�-��M�a^�\7��R%�=����
�û��a�`c�OĀA��ynx�a��/�9�7W_�8y���v��0�N�=�,����Ν����ƣ�i8N<Z�[�)����T>��`Jk�1e���5CPd=���YE�=��;�͏�L�!�f�z�2�;��,*�H��R<�0L�0Y<��"x������B��r�&v�څ�6���C8|�(�}�)>��3�ص/] ������x�p��B��8}�Ϝ��'p��!�;}G��3�p��M|�ѧ(n���rDV�����0<���*]yB��h�8��B������0��$�	V��U`ؘ>�
�U����^���V��IH�Z�A�X�>�Sq�&������%��r���	Y�����՘m2���导����^�K�[}h,<�u�/�EIU�k��W���B�e�SyH��Eee::�b��Q��m���݉.����1�s<�t�A�tM���Ͻ�	�g!��zBF64�����n���s1q�t����9�������>��-(nhAA���AAu+*�F��u<��� 1��	;O�C1�˂A^��m<�#�[D�������&U�m���54B!�:+��w�e�jM��Ʉ�^�pKj��~0���|�}0Y��ɇs.��! J�����G�7'��Uk���,]��t����_��]�����"<:a�x���J#����#��~�L���E���)*�����"-7[>ߎ�7�a�������O/��{�t�ll��־�8V/��Ջ���qX�`$^�݆ן���Yx��q���8�k3f�o���&�{k%V-_�y�'��� � ?҂}{����h뜁��i�Q�$����6 +E&x�7Yϕ��By�5���B0�]+O����?.{�D4`����:xF4SM������tep��oL#��3�	�s�T�� 0	��J�ܞ���^�]�"�@���=D��k��{��A0��k�ɖ3��w��A�� Q����a�=w<X��ѐ�Ėܲ���a�=߅a��\�m{�}����0�$˽�����7���-0����2l�����X�"܃C��_��kׁv4v>������6}��W����w!���;'c��#xy�0#����1��������h1��+�9�y�X��z�'����>

�1vL;���c<��R���s�ObђE�ю��Ƥ�Ӱ���ᓏ�:r���'��77;L���>�k,}�9�J���<D��!&!	1�ɘ5o����O��Nl�\tI��ja��*�!���'4�i�U[���P=��:6UИoGR�$�̓�5ܲ'��J���}8�B�So��]I��@�M|>\�_Bi�
q�+w��%?��������/*�����y�w>���"����ᄡ3�4t��0U#����*�OV�w��0,!�HҟQ'I�f�4he�zգ�N�s�xy�µ�!��@���*%���UOGh�8�Ĕc踹8p�N�����I�����ho���,�B}M=��Q]^��"��0m�m��=�=�"�M��ΎnD��#�+-�m8��8��,_�9up6���NA�5$qT�#��G0��x�j��d ���k"�lBYf"�ݢr�NP�{�%�bj�A�ю��q�S�0��j��؅�_�����앫��b�����<~�������c��ر�sl��C�9����i;sX����q��i�ٳG����뷰e�'(���%�Q����1� ������|aX:pN�������h������]��J�G7�^	��0\MΑ\�V�pt��oU��U0� !,?�+��C2� �u6�a�,��5g�!0&��	}tbS`�JBV~L�H46��0؁]{x���@{hu&�'�!%#)��HN�Dbr�������uFA�G�_ |��i� (����`��<1��������ЙC��'�� �>��sr���;�����͋򆋻/�=���� =��fxY�`���Q�+;z���	���a�`��n�1p�Dc��v�0$��,��+,^��&�>�Q�B�ː^3�YI�ٙ�F`�Q �/�;��X Ώ��+"�Y�w��?�a��	�:>C�p�^�q$�:�������2B�g$���A~�H.jƞ�7��ϑSъ��|�"R�1E#9���J%��3��Uj��/�ҵ�>DzA1���|v���<w
����T�	�%X��#\�y���ALr"f�{�^x���<v}������b��2��Z�5SK�Bg���'&����������+1jH)r�"Q�����`��D�9���8��a�CFO�Úd���;�������m4jGZa8���݅���ce7�L�p�˰��	�֩?�8���p0���X�<ŃĢ��2�^Q�0f��������|^��� ��?��?�~�L�<��&۠�W2���}0�&�`y�'���ʞ��	E���J��/Y� ���d{�ϽWn���a�� cLC���@p��0 S�ۜۻN͏��ZC 4��
�����U!�v�� ��'��{`��kݯ �J����c?+{�ޔO�ʏ����9��O|���>>q
�~�=�/O��-���EK�E��m�$\��Wl�b7�+�[�W܌`c���0g�Sؽ��^V���4�d4K�.!>Ͻ�6�L�}�$&D���?X��+W`Ŋ�8|�l��e(f�K�/G��N�陀Қ
tM�e�-���=&M���b��YH�d�m������p��c�̹�3|�����p9��s�O*g�QOn�%���a��k�K(ۗ�j8���a}�)0v\�Nle?҉��)�fv�'e<(��pN��S�I ئ�p�W�\��k�����{���E2/�����a��٭�Lo��0<n�,<��*,\�?�g	��[=��A�~�v�Z�n޼�$@l��S̰��_~�Σ�1��g_c��!3'*������W�z0�k%0����S����0�{0l�C�uW�R�6�	.K���N���Z��p��E�����j1u������ v~�%�~���PY.�:�k����c��d���p��U�Y�
�Ki�ð�8q�"n�`��G��#�E�<ʡM�R��O�#~j'i��R�Dl�L��#j��Yf�_�0ӓ	���æ�q��CJ��2�!��F�sh1��M�ӫ���gp�Ώ8B+l��}��$:sO��cp��A�<�N~��7��̕�8z�$�:��GO���;�r��~o��!46��VD4�g~�k'B_Ff�j��[;�.���8F4���Á�� �av���h�����V����g�L ���0<� l�W`؇e&og�!�T0Q���1�I�($�������RT���$NKPX\���x�Cà�!����#X�G��@�5BO�f�M�(#��FBM\�y�W��F*::����M�8�110EEB
�Ԇ@,�0!�hQ�Qzc(tz3B��"���R��Л�afGeM�r<��#��g��g�}	��8sy���>Ђ��9Op�'��5)�X&)�$B�%	��Dx�&S)�6�@W���zpMN�U��� Oʋ`�F�#�)Vn�a	c��'��d���å�%jt86 #�q^_	��8$�7b׉��{�J� ���k�V�E��aЇ�b��Y8r�,�\���>َ#'N��݂�Z�[1���@�up&��z�%)�b�����p��e�{�q4��^Y���.��%�e�X��9<1y(w�ᕩ�xsJ!^�L�ks����"��S���W���s�^�����V!"2���		��+z҆#�O��s:fh��d��p ���~0l�mEhq�hN��gO OT#\��}�=2Lr����.����w�8j���>9�7�=�Ai�Z8���F ��OA!ʟ@@pș� 8@D`�#�*��"Y��8�v�H6�A��p�&"�R.�NB�M���-˺]�}�(W�s�a�= ,�bܣð��^	�*��λg��F8�!��
�<&��
�V��òN)�~�5������?K�����?A�%21��x�q��/��l�w'��	W	W�ANu��0�ɧq��l�u Y%��	�%*]��`��m�z��8}/��!�r'!0�
�yC�nU#4�Ͻ��`^}m5"�ͨ�����k���g�p��رs�?���J�Ꚉ)�<���4���{�dL�5�<�ᙳ&��/>ŜG�#*.�-��=������FL�2���acJ̙�����C��&~5p����
�����v��{�F@��6%}۬Qp�m�[�px��V9��)� �{%�6��H�$� ئ��p�U��@���Ŀ�,���V���;i�,[�
O>�ì/��0,�$$L�ί?a���eH���f���� ��
�6��K�U8D9��B'�	���*0��m�bՃ!�&K�l����pm��B�oL���Ç�P'0|��������wc�W_�򅋸Dݺv������W�&?wn|�c��͟��ɋxq�
D�%���m��gn�[��k�݆��VXr���Mb<��U؄wx�#K_/�0,W?1�y�,#�Gx���LC�x��'#���� bJ������>�q=�-g�Ih�f"rk0�闰e�1������_�������=���3n��#���78~�".ܾ�B,.�ȿ�x�W��w�yE�m�J,@zq����%<e�j��Xa\�k�Q}4��U�q�ld�T	G�߅a��Vr�f�&g��K,����!
���CYfyp/��9�FH�FLDNe��2�㯁��#4��Q��伃���Z�Z-aa��_�U��`M&��H��#�V� ج���3P!\/����WC+k������/���뇀@�� �,<W�AZ���%�0�XgH��E�����(���`��g\�UL�G�^Z���.�;��������a�Kr6	�OC�I��H/D@x"����AЄ��C���,n[�2P��U�1�2A#� �,/r*1�i��̈́]��!���cǐ�v8�����0��`���}c+�Q�`]@r����������Q3�jR��Qp	4��'5�c��';��2�Y���ڏ���G�bي��>��-Ȩ��ʡ�N.�{R1�������_������'���c�֭xz�R,[�>߶	�nz//���j�Ҵz�2������rLo�ƆU�����x{�Sho-GcS1�Fа5��'�a�4p�:�r��5�<q�����d����7�� L�~.	��*/���ӛ�v�w) ��J�Q��b���A�T�5v�>��{5~��D0!�����t4a?���J� ��/"P�a��z�ް�y}�����Z�Hns�3aϙ�j��W�[��@���+�>����Ȕ3�W�[	�D�T0L�n��@���6��������	�
`�yl©k&���=��K�|�7�$�|��=�2
�����^(�%��D 1�o|�	���	Ϯ|�&���_��?a�p��40�|��O���7��=Ǒ�]�Ј$tO����O��ճ�`�&��%��O���9(���TLY�x���I�X��Z��$����7m���oPoc��#xl���PL��8�.\�q�A��	h6�gLţ�ga��?a��)8~�8�O�AAI	RR���qh+}b�ץwax�K�Ȅox�cJ؎TR|g"*�V����t�l�0�&����1>^��L�G��a���H�w� ����7`��d�b����坰��10�v�M�q�� �x���g_}O>�,6~�������&�:��ܹ�	�?���g�9~
=O<�`8Q`�yZ/[�cV0L���m0+p�o��>E���q��.��5՚x���}a�J�P]����ÛP6d�l>tٙ�7X��ax�رصc'n]�������'��-��淸}�F���q���_�:���X���F贡h%_:w7����������h�DZm'Bs�L�N��6��\	]B��{`�^��>Q���XN%&!�֦ �e$i֢YZ6�a�=��o�-�"�f��Q8��)�3�,ymVo܉���Ū�����/�ާ��e�l�}l�u [���N����'��u(��.���
��#�V_h�h�ձ�J;Y�����)�w����{a؛�taX<Õ�a�@��MCi��``}�$�����l��jd.o�� ��Eڴd��Y粑+�C���Y�3�Z���d�ǥBo���7��걘 4�듋b��iHLI&�*��L{�		��
		�N��^O�4�? >�^�!� ����8
�?a�G�	���� v@��$�f���u!H�:X�%װ���z��A2 ���d$���z��0��與;���\<�;|f$���P�Y.#�" 4�Z��"��Be��i�@}�h��s1}�BttNEvq#���9��?J�byרm/�7AM`ط�	m
�my�k�G�0	1V������x�%*�޿�Y`L.�����k�`撕0$�փ�kI��'�Ç;����op��w8v�[\��W\��g\��'�����[�PP���px��" �
ڼ!p7� 26��O�9�%˞Ų^Ħ�>��`����`�����*<��d,�iƳ3Z�|V�_��zZ���v|�n%N~�o���Z�QP����b�1��/���`�	��Q�8}�&N��#��^��z��x�6�e&��`8�
�
�{�$�������!E=�#����/W ���'�	��@+�bY<Ɂ�]S0�0=���th
��i*�
����|a�ْkUr�ߕ�қ��v�E����  ��
�����B��[0��3l���`��E�'�cW�J�Ys��$X��uT�`�� �!��k��3�� �<�R/;�y�	�
B���r��;��"����6���HH-Tq�������Q4���q��x��5(-mFZZ1::zp��Oط�42��E��}��9�)�&�c��1��#0��U�l ��r��G ե��I���7�~������K/���}��y����SO/GzV	
˛��9K^z�zE���Y��3���s��=��`ᒧP]_���&tO�Lcs$2s0�k"!�!�����ǘ��~Q��r�M��!N&�+�R8��1 ��0\��65PHp.A� H�%�p�G��J�d	��H+��`�{�C��ð���>��t?��/�v�8a��?
��]�'�}ϮY��/<���>��qV�
�.�ϓ���ð,�ا;w�m"{���°,��⚧#��
ñ��Q���p6V����#�ˠ4z.�	����� ˠ<7AV�������f���m%4bL�ʾz������Д����Iط�(�>��	�W/� �`�|�=y
��ȿ�����3*��7��÷.����|8�oQ�q��M����h��nŵKw��zv�S�T�s6;��z��H|l���]��݃ax*5��f>��H(b�T<�n��g"�2p>�j�lL#K�#���'�Q��S6ђq"g4BR��Х6�7���%�-GH2A���ӈ��F�gת|��� :g("	��ѵ�$�">o,RK& �b2�+� ���o�pv�#���^LT1Á���5ڂnU����3Xa��^MC�%��h�+ϰ�N��ñ�#Uޭ`؇e$���)�/`�9���BU������0c�2���&>zo��.�o����]�����v+W����,x����`0��t�+l��`�6H� ?�7[i	�^�B'���`�l)�p[�p����!z��=�}��,PL �p0�\+b}T2p���pl��F�[���C���h��N�m�h,]�>��_8���.�͛0jr�J����'�-Û�������ٗV`��e8x�>���n���[����0y�І��9(B�_L9�XW����P	��p*�dB���+4)�~�`8k8C����>�Q��c��^�<N>a9����]�����'�����VF9&.x��}G��kt�{cg-�����������%\�ز� ���u���\�p4eB�ь�����EQI>�t;���]�x	چ����s1aB7Fu�a��x���̓�����X<k^]2Kf����c��.<��\l۲m}�=mhY�gV>��-E��Q0���c�x=z���t��i��(�����@����U�:�=���w������m��R��@6���5yS �\B��?	>|��	�^��=sƩi���[7�	�֬�TZ���	���xno�N�_��M���T�&�q'�/a�#��{����ma}0�e�ɿ&�J	h>��]�(�����+g߉ ��kq�u�)�t� ,r!����Z2'�-c��*c����C� 1�
W6ؒe��O����W$�a��:
n�t�f�a�G;@��@9��u4f�Y� �����S,X��M{g����]�0|�$̜���^×w��UOcH�0�M����_a��+2m)�� ��\�r+�j��j`���lEfz
�0fT'Z�v`\�T|��c̜� �Qi�	
G�)	�|���i�>	�I����g5��/w`�o�i��9�վ��>�D�ģu���rg�Xa؟�|@�I2���{�Jh�/�`��婆}a���R:������/_�����JK���$�
�zD+�3�{���m��@�w6��7+�$��waxȽ1���?Ͽ�/��m�a�_ąs�H��&��[��0����ӘDN�������?����@��]	����J�^骨�Y!���	�F��m(�W�!��@�0|WͶ�$����d�Е� `ς�p<<"�Q���G�c҄	��°?�|�1�<zW.^ĩǱ�����_����y�:n\������S7p��qܺ�v~�]c&a��Gp�·��;�Ϗ �xv���ψ<D���ɵp3e 
WC�/L�0,�E��B��0�K��D|3�!�����e_81U�`ΟJ��1�Ng�:�0<������*�����Hdy�e䪘&���!�a���1�/�Db�8ĕ�B�%�p4�2�[�xdT�A^��V�N䌇�Vs�x��G�P:)�%��\E���E8l242 ����ĆV�O<�1��a���+ƫ�ck�[�bOm��~���4��ap1�A��E�7�č_���/�Ć����^~���ؿ?ߏ;8}�_�s���vT�����:��b�Gf�]�wa؟�#�a�x�M۔�dĳS0r[?���x����yx(�6[Ba	CXD�c�`" �����ZB��
�6Y�i	��<|�	��j?�� 6��|��?}���Ե�}� ��*[�����ǀ�<��K�⫝����6b8&����e�j0y�4|��.|��v$eU��7�4����Q��QJ��a�c��6���j�;���Q�P�B��`8����aH-��u_��+��]�?�|v�/���>?���s����~�ͬ�����q���4�GN���!(��Q�.��L�!��%�ؼ�c\�q�`0Q1�O�t��hl��S��a���1{�XL�nǔ���،ntk��ٳ�9�����r�x��W1n�HL���|�����k�[���qSs;.��O��N��b΄Ot1�	��dB�߀a��J��	��Á�Y�O�ȟo����wԝ �o�7ʓƨg�6��Kx��~�j�M���i.��!�9u'�)��U���)��J���Nyp���o	@�mr�\y��)�O�c�
�E��Jy��a�9�a�X[+�:��~�F�njB�x�y�<�U���VeO"��'��Q�NH���$�a�w�~�B�߂�q�hY�BXs��N�����ym~,o¸w�(��ݜ��S�q�.~�|u�um(����.�����C'�`�קpC ��M���gؾ��_��O��'�Ɖo��̏?(�����#s�t8%�É0Uބ�?�\��m���3���	�����q���:�%f��+v�Zp��9 ��1���V	_�`�{!/3'����3����g���m�َ��e��O?��apf;�Y°�QT'3ߝ�:x���h��{����ԋ0�-��ic{R�b���?����W��`����a�~�+��r8�/��IɶA8�.�x���p��3���;w�Y�
�x�Yl��c�&�t���	�9�����&�V0�����u�{axax.a�Q°�I����E�����k`�� <z�nV=��GÜR��9V0&)3�%����lb�l�~�$װ�(^f�<fa7a�5�����c�=�a�X|���G	Çp��)>��v�ıCp��E�D�������~�~�/?��-�>���v�5��]�p�����N��M_�l�h�K�b�`݈�!S[<��2B���px�LñM�`�e�2t�ǽ�V��6Z�Q6���#ɘ��ƧS>~�c�S	�S8%D��@x�LD�DHz��Gs}7"�&��N4�x"���#�d�b�I
s�hD��L�����i�k������g�������ÞD��U�#�ظ��;c�
��8pm�D�Y9G7�1��QU<��p%4q�0�&j�{?�'Dŗ�	��`8�ѽ�nx��������܀��i0d�<�M��S�m®�7��q^{�=�5s�H��|��w8'/�����/PZ^??�C-�Cl���|�IB&���`4���@(�t�@TT���PT\���$��B������i|B�s�PRZ���<�A�/  �����~�R°� x��	��~�j�0��>݌O��=��cö�:�	��J��)�m �Z[��W��Íh҄����z#��`Vf66}���AM�(xhc�O(Q��|�J	�e�N��_*A.��P\��Fօ�0		��s3�`8L��������hv��1�.���T��%�"0���D�Ɉ-iŌg� �����۟"����j8�1HcF[�v�����G�~)��+9C��AÊ]�x�#S`�1�[X��֭WC.�{t�5pqsezAoBvv�Ӣ�����=�AC(Їƌ/;n�`h�K>�~�%�0dL>� �GC��cX�h6���ax��p2��+��퀌�HB��$�8�h����*�J
aX�$��)
���hqB��y�D�).Sn|���n1n�V0.y�:B��%��I�o�V�r[�z����V�J�u%���[���Ly|Bb��x����wș@�D�s�9�	y"�ީmޅP�J ��q{�g��Uj	�V��#��1��O"B��ɑ�8r_'�Y��c;g �4N�g��Ʉ�IpH�WN�)��z�zej8��]J���r�a'°�H�v�l@�J8��9��2��}���	�>i�4NG�X8Ӗ����a��K���t=���C1�Gwc��xo�WX�c>?v	�2ݴ�0^��9y�5���3�ᕏ�aۉKxu��M}!�#��Z	Ǹ\��5`ٛ���ɓ����hg["!d^��pv󆝣'ٻ���n>����UG��E`D>ۖv�;��ps�\ao��Asx8�cb�S�ҙB1s����N�o��d³�K�w$��"���e4���n�&e$4ߠ̱,�N�r�NNON=ه	�`�ސ��t����X ئ�?X�{���C�U��J|7�D(V�@6��54�&�xNb���;0(i�=����51k:��2�?�4�m݂�.����8K��������l�?����F��'|}�,z,C*a8�0�4d&��EB�|��#�"�Ys� �XZ)C)O#K,�d8����x�o�a�|�ջ�=���]o<�����ma��RB��f���z.t����x�MaK� ��;�_�a�u��d�S<�
�+	�E�ױ�}*��'��Ĵ)��&�O<��ڏgO��׻�o��zN?�K�������o��?��7w���]X��j̛�8*h	m�������_�n�n�6u��+�\1��:�QO��lT#�HL�d��"d�+�P0,9��i@�A��e�޺UWC#�e8�ޔ��������Q��|L������z�ܩ�k�ٍ`B�kD�"[��l`C�c�g�[>��q����6�a��v���,;��I�����Ir�v|&A�;�9�xPh5칯&O���l��}d-[$�,a�H Ұ�I����3�OkV%�r�#�l�
w�X`I�ft��e3By���~֤6#�^�\-ХTc��5X�f[�
V��>&M����",_��5h_F�!�:skׯCIy$N8���>�� �� ����7�͈��Gtt�c� ��)))���D#��z�A�x�5��.�&���(-+Q�D����70|w>D��s��\^W�z����xk�;�}d?>ۻC�;�CUK��㐚����\��<O>��֬����ׯ��4�=�C[	�3�`��۱n�6T6���9����f#P��IU�J�z���3�Jc�p��(!0�)ό�1���S�d�(��pa���Q����Y}@W�bh��#R��%���&�apH|	�q%�4Ɔp�|��SX�����ڄ˄���i�AN�Dy]&�W5B� �3G �pͺmJ)CZ~^�]\f�����ȥ��AC )#�qQH�LFt|$�f�}<���I�C_��11�|��*m���7tQ&h��QG�[����4B͈KL�cO,����q��e5�� ^�kx>;�*�P�~�U��U4줬�h,tXc�ՠUpc����N2٩�=ʙ�@* �G�IH؃x|��.��]����^mrV˄/ʵ���w�U`8�p'�K�tΓeBj��U2�B��S�A���S)��A��
P �e��h.6��\��&�~�{�q_����/�R���;o�M+pl	������!{�EY�`��	;v�vlOE�J܎+r��1�ח`ۧIpL'|��z`�.�ا��bC`��Z�5A������^AJ�H�9��S�{�b��׃����|8��u�\�����#��#�m��&���p��e[?>��J.GF�x����n�W���%�����a�9	��;h,	��f8���)h�cB>�d[�&N������G�~�W�~�_}ϭX�%ϯ¢g^Ʋ��`�k0��W��'^���0$�- ZC�vM��I�0u�,<��i,Z�K_X��o .@ѿ��w�o������.\��3N^�	�]bۥ�K2�e��|oZ�1�|����R>�'!�Ci��|0gU'ܨ?�ـ��߳�����"^C��kB��{���}�W6���:�X9
�f���$ �����|<j���a�A��{`X�W��S�p�r�yj���!�^��<�gΜ�°
��w��a���4�1���
�6������W���������3H���pvǣ�GԨg��]'0<� 6�����U��S�T�0#�ф�H����T�cQ7���D�l�M�.fA�\4�/�tDU�A8� l*%�r9�v>̵�s	³�%8��{�� &K�1ɲ�+�q/���&A��%g�.�ͣf� a���3�5� G�fL�Ɩ�k��0�����ҋ����hi�{�l݌cGv/ ����n�l��G�ä��Q]Մ��&���m����{Q8���MH����q��[�a��y`Li?��y9�~:b�g"�f���,�Y�ȻU�$��a`��4
Vv	���O'��_5��K��=;�v�<B;�A�
�E[M�(Xd;�jD�d��@�FH	�Q_���%$��!��ԜG�Mg��rb9]0�b�b*`g�u�c��JY���^W��B ���ͳ��-%*�A80��DaX�&K,� qhn;bJų-#б�e��s{a8�_Rwɐ���	�6��[|�x�G�=�&%m��:~G�~���#����[�m�>ő�G�㫝x����>Le�p�Q�~�}�l��P>!�i�,�%�!�}`I�5[,�h������q����@l0���T������*�IPP���+�!�Xb�L�P^K8�	�A�4Bx0��_R�g_~�}�������s�u� �������a�h;o�}/�z3����5�ⳝ;���A5f��O=MH~��y�:'���7vX���M(�O�U`X��|�&A �%����0����j��&0\��0��K/�w�)���L%��D�xsW���:��sh�.�5��G`�&E�N�e}��NbSN�M�@����?�%��+#`���%�'��=���)|�x�����\��&N_���O����㓯v`�_b���X����a�߼s.���� ��%Cc�g@�O����x�o��>�F�c>ܾMپc�~|��^=ulrq��E횋��4D��'Xc- L�P�&���\{'��=)�}X9<�y�Ch4��=�^)4L�I�N�/%����^�`���j��K>A��, l�aB� o��>�Q�lG���5����L�a9{2�il�gM��L�,��� ��� �6o[��"9�[�b9���B��Y���煵§��U"�*v�`� �$�6uSa�Y`��v�,r��5gL!L!(���=�����<���<��q`+;e,x޻@,^7�^op:��Ra2M�1C���&�=���J��n�o�'��I��HO<
.�mӈ5����;!% �!��ؖۙk�*���2��1���-4��������LmÀHn��ka=�oC`y;��.����Y|q�6� 8���8�����ݯ�|���U��ܦ�nފ��?�������X�߃������Ϊ1?Q����"����o�Ǖo�~ĵ����i2��'d��x4�y������O�[���	p
�Y&R.n".�n�����^�޿�$�a�^g^�u$<O}�u�`[2�5��hJ2��XOz�iM(P,�b�_��;��dL��w!�&I5�G�f}�,0�r�9O�^�����[>�%���?-�b���.]�����X@Xܰ��M�&���;��o:u^�pz�X�6O��-s	ó�3a�Q5E)�r2�w
"	7��S[31�S	Ta)�$t�&(Y�4�MJ8k�'�5�^$6"8��b'���B�?�G��C���iw� �@�|<7���ДN�^ �`h&[�V�P0�!��e�9��-��rW\g���*`צ��a�t��s��z��C`��a��z,|t6�zb�̜���c�G�|�2���J�޵��n�!mX�� <c�ta挹���GNv	Ν����~�{��BJ�ph��J/�κ>�/YB��IT����1�3�2���C0�K�T�I�D9	�=JA|	L�S��T���bG��H�X2���v&Q�p'X�1��LT�� q�:��;a(<b�	0c�<'�؝|��Rv�B�7�m��a��`���!��lX|���	楼�">/n�ǆH`X��]a%���\NH����x�����$�AK�Ii 7��!�D�8�Z4�|��*X����j��^��a��b�u-�ېZ:q��0�'������Gyy%F��9�<��ӧ���	�	�*�@>����L%�|�&�]�W�X�u�U��"�9X`�PI����RP-����a�_�����}t���@vN&JKK�R$%%)6�����<~��4[������Wwx��"".�g��3/-���cO/Am[+b�������VV"���\�,�>�LŸ��PY����_^���zD�����l>�2��x�+��+�b�$����0aO�OH6����V�(U��X0�0\�H��(��ϗƍ:�Z������2,��8����#���H~ޔ�n���\�Gլ'mjh)O>̓��<bjx�
ؙ��<V|B�KJƢU�� �7n���oq������ىKf���������?�8���b8���5��7����d����C�Ɖ+�q��M����X�n���[����o�y ��f�N�Ϩ2�AuZ�e��aMf�,/ߔF���h��%���m�{t#\c8���M�՗�O��r�]����H�KP.�ݕ��]	8���*6���6�&��i� {�E��W�xs�7!ٻ`:|(_�O��i�m
�# Kx�"�~�j�"�J�e��K�}����A\6��%B��'lJz2[�
O²��;w
��dރ���	�&A(��N���a�{�\'��5�p�$�0I�V˽y�؞4D^j�r�� e�Kc�e��s�\��܏3�k�2�/��3s�ye�̶�9�p��#rc[��k�}��A����:�^��Q>4:|h���=	���O°��aa�g�8n'���q]5��/�W:�rm�D��_�d� ։@�wP�D��)��k�hJi��ؙ��K:�}�W~KeĶ�E#}���c���I|p�>��">�s[����^}��6|E��V��W"(���x����M�S+_ǧ�ዯ�`�c��җ_��_���g����X��N4Nx���i�������k"��~�)72���$'i��[%�P�^��{`�?@��f��O�@��{H��e��d��:�4�'܍�k�p��0u�m�v�pNJ�r+�=n�Y�n+Ƃ��Se�������K˷?��gx��%Lb�,yu%f-zo�/_���d>%�&�G��/?�����g.`a8�q\'}�-� �q�-��Y5���]=᥄!��
�@vB��[�6�q�в�N�Tq��T�c穗N��Oj����&���&��p²;�?�E]/��0`���/�e/�Wdas���	��'��l�F����0\!��`(��k�Gu�d��yPy���3��Q���qC1{J7�7˞~O>>O-&��ּ�
���_���cƢ��55�(�/Ơ�N��MS���~U���s���Ɏ�e�Z��"v�e,�*'V�@(Բ�����cf"���A�LD�Ρ�@」�6k<����L�t4�ܖ�+1Ě�n���BX�5�z��)��C��� ���5��u�8�L¯�ִ��Gx9n/�5�,����
v�B��pKm�8n�M��	*~�T4Ie��r]�dgma��E��ñ�a��A����>�g88Y`X<�V6�r	��QN��aaJ�ړ �T���O�aؓ0@�N(�>>��t�C����NgBRb2���QV^���
d��`����h6!�0+^`�_�Zc�Gt�1�J�(B��m�H�x~�##��HJIQ1�ń]Y�KLP!�Y�h����^G"223K
��Y���,�>Vy����0�9�+ �do��F\|��3��2�7Ak�/������|�$�AcU� S�-1�6��͔����]�d=�`}yRVϰ5L�Q�/��0�yvT�Y2 ��yVve�U�(�px,��iPZ#ۓx�k�%�5LD|�X8��^`��0�z��{}\-ENo�!8����6�d��r�[�0H_;C��#��I�E!F�}K�X���݌�k?ƫ���[��K�}��ي���Ս_��/c���ʄ�9Qi���fL�y�^�	�l�olڎW�n��6���'X����q��Ͽ�]�#��.�5Џ܃�Y�.˨Xl�>���]�Mn&���5��e�Ȳ��sL=ܒ��3}8ax4At,a�������	���|�������	56y�����A�Q�E��^/����^2�!X���aO�K��#�����q2|��c<���`�\	Y��T��/+�Z��cy��cچf����`��-���w���w?w�_���ݬ��b�Vɀ��&����bW��uٗǠ�ܒu�3���E0�dYe��VY=���	���*g1�_�|,������HuJ�L��=(�6�P�|N<��}��l)��IC@�����I�&{�=�W��܎��g�@����y�^/�x�5O5���ō�������y���z��J���5k$�Yל҆�9�%�$�	C+u,i�Oa���P��8�;�@I�|���UӢ���B�>�P�^�m0p��f��_����j5�AY�hT����hՍ��Ѩ�r�б�6գg!�u�v�C20�+!������Yn��,Y��|�֡�����B�M��| �!(�<����@�I%����a�u�p	��|x/��'�t>��vx&H�	�����0�
/��p��l##�����1�
��G=RZ�Vx�=Sy�M'�
P��#��y;evи�Ne��{`���6�mF;�i0I������ax��'��B���Y`X�I����0��O?���^n��~0��2��Wx�Rd�D���1���[
��\�E�3J(�%��9��ΫFxf)�)�0'�!,��TQU�ȴ2D�W!"��9��I�0�C0�c�dADAbʻS5Q�5����z�@,l���d�,T(�+� Z%<A���S���3L.��b\�bjQ9d��a���g�ch�N���K����`ͪ�a��x�x��UX��M������*���¼|�*���KD�����	�1�|ȷT6�w7�Dx;3s:;�
v���� �e9!Co�a&S7��W�S`��=J�-�@6�����ꂮ`
�e�`"������!��g��6o�
k	�M�X5���x� k�@�5��@W���hJ>c��)��;�:���m4l4�١J��LC�	��,O����e��#��*��s���:&y�W�7������� �a��N�ڄPZ�Qţ��O�0�Aw?��s*0l����1�oW^� ����B��X��l�!�F!<<�ѱHMM#��!:&Fyp��+@+�^�	���2�2Jp*��6��`�z�%-�S��a�����а0?Z�N0H��� ��!*:�qQ�����("���XZ��ҽ0,����y���C�����`�䂇;���?�O���<X?}�!���!46a���	)	�BDB*�(s$�I���G%"8*	����p	a�Bp��z��'Kj5��?{��	�B8�°s��������V��k~�jHgMZ�b* �3�W٩��?�'�N��γ	���{C.�d�C�6g��7���$7�)���U�1TF�*��1ޱl���"�b"�""o�
Z	�m0��+�� *�q��0H>p�Q��.����4��vA�ɇ&&��Ȯ�@|a#�
$=a5b9oN��'����Ef�ɘ��������{aX�6�s��8X��Y��2x�X�����F����3�#���N;���U�hj5�0;�%塼:�|_E^o�U�<�-���[�
���jJ �V�olSd{%�=ޙ<!Û��ũ'�ҝ`e�:��i`��x��6H���B�y����ݗ��#"�x�x�r����)��;w&a �*�>���r��]�!�ZD?�3;y�\��[�l��T^����cB<A��]J�����~�gr��c�
p*�u�(;x~B���J�p��Kj/9�@� ���!����<�g��B��" ���#�FQ�q�R:�Ny�^��|	�i��4�$l+�lO9ʵ��z	����{�6���l�.�Za���x�'��1{��"��x�c;=��Lh�ot3|(ߘ�ƶ���n�ߘ6���e�щ��|�;a���ME쟀�����6�i�$`���`�]PD�-,��lwR�(p�a]�+��"�U��ƺ�&F�
P�[<�6��oaX�g�0,lSٞ�?�Y/��G�)�Z'$�ٖ�B��n�4b���vB�^��� �|8���d��ќͶ0�L�����<��嬎�jx%�����N!Цu�,+WJ�Rgh$9�~<���ao+��3\���Ӱx�
�z�q��*�υ�0��/X���0���&%O~�d�ӛ&!�0�B�o��pT�4��$�V�(����ų[��}\��)�άF\Nr������XD$�#>=	T�LӨ�ħd".)�����|D�� :�Q�%�/�%�p�Z���fD�@|�x��OAT�t��C�f�	5waXq5!N�tLBX� pa��ש4kՏ �x��Hk�P;l��}�h����y�z�i|��G8y`7��;>݌��ŗ_l���6���V`���HIIB(�)��&QQ�	6b��@ť��ыj���BlQ3\B��#��T���?�`1D�S�52�@t�ܯ��a��h�4�J�BS �������?I%�W��	���S�-���Ѳ��?�ɟ�4�RM�x�ue=l � � ,�ZW��7\,#^�t��
!������Q�|N)�mv��l��I$2�S�@��*v|Q�"�N߇A�6B�R0L��A7�qÍ�HHD��l6����Y��0	'���0, ,
Ji�6�!�M�g4�0	-�.�u,���dBm�0�B����:� �Q�QÐ�J�:�r
K*5�[��$>X���C~��U^g��.""Be����P�'���U6��r�2�����855���cs�~͉��°,��0���G����3�<����	G7t$�;����ЇF %;Y�ňNN#'B�8,6��B8b�ҹ>	��$�D� (*�����°O��p=�l0��S�p­�a0g(��C��������W�eg|#���W͆��\��	n�7Ѡ�*��!|�G`@H���W��i�>���One�aǝو�.e�7�~�(%�@AdT5�#y�I��&$7��|����I�H�����o,׳}�6���+�b�{]6�	宖<�&�Q�
cF��%�u0���l�u)p$ ;	�&n�O����<�^|����������w��APf+Ӈ��X�>�n�5p����R���R��ӧq��vH^��Ɨ���'�,��>���& �Ժn,��K�qܞ�ĩ�,S>N�]���1�o�(u./N�8����J���Iy�!��	�2����'*�p��+i�|E�9�"_�xo�:(o^�\�M^�f%ާH<gV������SY�I��R���N�!�pٗ�G����Cy��(�PO��]��x,^�URV|F���x�z%����^�uJ�If=��|^_������y�x^��/!S�A�q'Ըp]������p�$�d	�pJ����+��n��]�΅��r[7��]���B8K�f���ɟ�4R�c�r�ʃy=A���TkH��P*�@}i\�gL�&{*�{B��"(y"�{����χsp:<	hA�H(�L��Ւψ,��E
�h4�J:�	��YGU\6:	��b�5���۩@�
����6��aX<�΄aǤQpL���&���uH	��p����.n!�T\�S�M����}2<�,G�M�p��s�8��?��x��SY�
�Q���s�lc|���p�! {���g}I%�a%0�6G�%W0�/�u(��a��Y֘�Y��{7�ƭ۸x���(q� |Q>d���0�4)���m0<�0�bg!�0l*놱���.Zr�S؈��JDf�"2��Ye��4*���lK*��8��;�b��N�yd
��̙=��=m��(/+E~n>2�r��@@��s	���σ)6f�qxfb��#�j<�� ��
�&!0l$ [�j�Hn*B%��b��檱0T��F�{�0�T6		�^?|&�q '����w�`�'�p��ܹt� �|�16}��~���^|�i,Z��z�HIHBTh8"�#	?� <��=B-�ػ�8~�X�e/��F�fG��χ_`���D7�L}D�S_I7�ӎ��I
�Ck��𐐲).��x�%Wr�j�Pb�+f�X9J��K�CC ��PTDl����	<a�7�h<t�h��H+"�j���
.�62/����	�!�%V�d���#�j64E�@7TN���Z-!�H�pyo�p��@K�@��&!��M��-KZ��0�Ko�l	�"%�Ot��0G��h! ��
(�f��S??�>�`��m0la������%�A�9!!���
�������LHEQq�򲐝����Bdd���	�Ζ9�w`Xc�aw/î���������\�0�������t�����`��FXL<���0�wXL���px�Bc4�3P��D�7,�Z���pa�� \��k��r/��#�B��,��������|�*��Ȼ@I�D|��4NFF�4D���{d	�A�0* ,�]2���=Y\#	ŔgB;�a<�H��Qv��*!�5��fv�#T|��ʇ�Nb�����������`)��h�����0�N�;B�ѱ��h�C�l8Z�#8��/��؊ш����N�y�,�(���B�E�ڋ��e��R^+����%�T�����@j3��x���Oʉ^��,7��f�� p'�x�ȟD�R�~����3���#��>^)#��5��r��O�i�&�&��}�y��g��3��ds?ʋ�M�Y����=��Hm���G>i��2m��M�-b��d[�_ބ5o>[ov�"/�f����*^��_
A1��O���+�p�B��U42(?��k[�:ޔ�(Mt�9�j��e��z�@�W}�D0��z��zR���'����mDr>��;Aۛ,�)X|	�>\��e/���=��y��D0v'丱,%~ԝ˲Γ�G>N��A0�J� 	�zt|��;��A��@*�F�6�p,�����..O�w�X�s'��-뭫��!Yp�g�SҮ%�"�j$�=�^�Jc7�m~1�_wR�����Y&V� �I�'��~!2
��)����r��i�dY���S�(�#eO7G��/C`g.�gH*|��M��&�1p��{`8\�-p�3�Co]��g0���px��k�6?~���͂wh.<Ë��d�D�Lh��
�S7�1	���ɃƉ3���{�$
k1r�l<�ƫ��d1�oތ[����+���.^���=�Fvc?n}q���Hv v���9��	�%���'�#��5�G�k�|,Z���<>��M?�	.��
����ӅS�q��gرm=6����_��ӧ���9��H�IB|lb�2��ȤB���!,�V}UQх�کb�s暙0�u�@*���u#��R�m�pB^;�q'��΃�T�k�0\�8�ۆ];vaݛ��}�z�߱��m�'���;k^���g���g��g8}�)���hokCvjB4H����d���t��g ֯�W/����~���|�٩�B�9D]+q�A)���*�����a���Q��{5�΀�l2	�!���Y��T
&�ڦ��ܮ� \:A���K&Q=$�ZE .%�VL����n�TNaM��'YE@�H8�}
�$�L[$�f΋�2�d�0�<-3$�x&�r^<���)�3<P���Ò��""1��F���0\���f$�ܣҬa	��Va�*N�b�(���f���5��M*sD�y��m0,��Dâ�t�8�{{{��lzC0��%L#Qy���3T�p|B��&�M��z�	�..npvv�����/������p (;I(��7��5�	ЪeSD$����������!*!q)IЅ�"�����p�K.��L�K*#��a�%�_]n+�}n�ˆ�a�v�������T&���F�V�'�<��\G�,A0���R�$�]�ߖtz~�O���,FW���o�� �5�.�up�%����!9���=�L��h:�%���w%k
�E�a)�/v؁����_�h�v⯺B6��*�L ��R�����t��'�P(��Dc@�����'�Yb��+��uRwUF�?ۀX$@ �2�9��ȅ�qc�&\?L��PW�=�.Q�Tﷁ���'�h��e�'1j�T�]���6�1�6����g.�)����l�:�����+�x�-G��S|����m��},���XI�_��1�*���>9�_$�15�����r�\{�}סd�>^{\��^�|%ϹM2f���ȹ�\���\�O��k���lr���ȑ�D�t�l�m�� �J�͑�US��&�Á�s��9��_�xn#�̩�ά�2�-+q[9��ښX�Mp��!O�IBe�j�5���\�S�N��)�Ή܎��cB+o�;�5��%��/�D�D�;�ͮl��dX���`���5y�2�#�m��i��D�cpp�B��lʂgd��j$ԎCpv6�c�%�Ϧ���2�4R�	�����>��9�	�=*�� �a��V ��;)uZ�9P6 V�oS.)ca�Ё1��-���F����E��G�6
*(R��M	j�������"�W"��iY�TB��1E#�� K,��Lq<�
�^
��Ѭ|f��4²G�;�W�&Ü��Ƣz�}|>^x�M<��l�hnݲ��9�
~��p��¢��U�S?}����>�8w	a�i-�	³�6�I$�>��������nFPV=y�+iBJv)�Ґ����#;���Ex��ױ����ܼ��/���7��[�q����o๏�����;��ݍC8yh6�O�\:�Z[����psA"�iňJ*�9���J���S?��3� y�%o�4�}�n �WOFT�x賆"�~��y�b��DD�D�t�x�\�O!(5 ��	�ݏ`��Ǳ`��x���Ɗg�����g`�����3�����˱m�k��W0g�xԕЂ��F�6��~�-���h�!æa��bܬ�S>a�4#�:^2V ��.�����?"0�J}����B=$L"\��u�\!p;�S(MaW$�X2��6M�z�d�@�ԣ$��-���'p?�,AU���[���l
���"���C�^b�-U��ɟ���)�v*�	h}��h/gGRo?�����+B��nBs�U|7��߆��P	Cb�%��a�@#���嘾p9
k�0l��݅!-��8a"��g��/�駗`Μ�>���*n�b��d �%��[�[� <"Le��^�Cjj�P#==������4�������ch	���e!#=��El5*��<�N�']�^�VC0�4����O�����npppd��	�)i�mlF����Ս�S�����z=<|��6r8Y03�����3�`�<��y,e9[��|�tΜ���<8�	����'\�t�a�~�a_3"].a���;-�H�P`�p����^b�G$���(G	�!$I�a>oMz$_q@J�%�-.���e����h.��"�>8}(�4=�sE0�������6j�_�s?Ly�Y4��ǫ�nh$�(O������i�����9�`�ٍ���eѸ.��æR0���R W�7�[���X�	}�8dW����o�x���?��<�n�Ğ�Oo��r#ˁ���FI1$$��cO��rvbY8�V���"�E\�(�C��E��);K����w����}Y>���u\��P�X�c�4��F�a �܇C	��$��Ra\��"@�)��B}�J`g�x}v�_M����c�ٮ?���V����ʩ
����P��YD�h�� �*2Ua���R��ys�,����qjg��99e��K�p^�Ʈ��l��e.�}*y-�κ�]�E�1Dr=�`*�U�W�]�����=d.�_��X����s�cP�D<�@��@��0����T����}�BC�!�xWY�<���1���E-�"j���yM<�Hʌ�<���^���|��"�y�j^�%���͑��v�Hγ^��}���`��/ߋ�>H՝*���4����/��!���˂3�u?����!�'G�������1�eR�?��}�~���h'q�_'�S��m��"�����Vд���W?&tZ��R��|��]��{� ����������r=r\�PN�p"5@��S�Xfn�� 4D��E��Yhoj����x�\��l1^[��zc���[o���/-��s1g�D�����2d��"",�}E��$��g(ǒ[D�J�h ����E��pL#��=u/����O^;|���1f�<<���x��g�A`��7
�%���0lS�W���7��2�~��cg.b�#OYax�D�MFB��nz��	l�[�ͭa'Wc^br	�qih,����`�֍�}�0��.~�ۗ>Ƿ�����M�ua���1n�݌��6�u�܇�~a3n_����?~�?���\�7.�7v-��5����N�FjR.�
�PS\1�/���I�k��¯5n��X=q\�.�xv�O.]�O���]��c�+��f8J���7^�y=O>���V�)0�$��t�]��<�U�����ga틏��ᓗ�ೕ�`ǚ����g�ѪŘ5z�i4!���n��Qxhp(���F:"w}
5�<��V�]���հS�'@h��i���Wr[��L�AF�U����`X˩����Y����=*݅]-�C[. -^cY�ڻ��\G�V�������@��$k%>Y��%F��I��{��d�LS�r��� 2���ś�����DPB5K�ѱ�ק���#�x,a����> N�A8��p����Հ׷����W���7���ص� !�Y��r%.]8ϗR^��8u��b���ʀ����-]��JȐ��������D!!1y�9
v-�T��ظh���=�r1���݀ �tzB9��D*"̄���&'����Ъ	�twE ��T>��/a؍�����;][_�U�_��={q��I�ڷ_�݇��wat�(������w�������xo��x��ǰa������xq��xn�r���ft͛s�M��8���'��R{�Y��ѕ�=�.wA�L���wp�BI�72��[l���Α0�&0Ly�9zK�C��|%�X�+�ZΡg�"@�,�XE�4v��+��:�%N�'Ir\�侍p&LI�q�,Q!�)-б�.��|FewC2xKf�l��l�ةz�S���/{����:K\#�y�FX�Nk����d�Eǘ:vX��*xH���2%w���}��>��2�b�dRaPb$ȇ�|w�b�qgǑ��D q"�9p�L\G�r�#aÑP��6ȉ )�3%S�>�z	��^�T����羃	�";��h�j ��a��C�"U���P��Nx�B�Gr([%�v
�)�?����v�b%{B�=aN�6(���C������;�l"�.6팄S#�����	��,7{��eϲT�Ω ��P�[ �Z�����M�Q�X'�1b��t���m9��;� :��������Z���s�(�9�5�eى���H��j, ��g}>A� .��!|6!|&��Az������@�zHOq�������>�?�|�(�+Al ���)����|�%�����)�;^��{;�����L�=�Q���\�����0�p���S�{����������f�"i�$d���aW��.�p���,�}^aa�-�`�'9���C��(�F)9fZ�-]b�	�i#��yg�Yp�$�#$����Ն!D��8��g��#���'����8���8�k=��� '�m���q��&��߀C�����w���W��ͥX��T���b|(<�P�>����T��d������#��D`O�c����
玆]Z���0<>�C��?K__�ǟY�u�ȁ�n*�x������`���a�6a��M��O�3�=g���t�p!�\)�# ܎��z�V�"�����c�R�>t־�� ��׎�K�p���zzn����o��G������vB�v5��V\9���ܺ���܁�o}�n��7�w.�������9tr2����X	�H,�%���zD�@l],�ULmd��4�FT�6�*��=��?�=����� �����KVbȨ.�^��܎/�F��G��% �/E�5�1�O����GF��#�ܜ�xq�(�0�/������C�hBr��� �{��C>`���'���s@����C����
�z�Dj�
� ���T|�`�� 0\�{(V��̆�z6t�3R>�Om�S�U���_�ߴk�4�*��@��r߾�6�Fm� �˽
pmR0la�^Y�mt�Ө�J!�
���8������ٙK>�7Hr�&��#TH���p��'Mj#��S)��,�gx�ހ�W���m_a��S8s�V�X��{gN�ĕ�b��Ǒ���fͫHMK&`z�l1*���šۤ���dbb�
o(��3#D�ETt��c��d6�c%%��cx�`«������&�FC0
rPZR�(Z�]4�����Ć.��2S&noDP��^>
�%7��pGG��ۇ~�	׮��񓧰uۧX��)$������1�x��yx��5���mxg��k�BmS�T�a@i}�Y�
o�)�ɰDW�'�����0L��a���峐�f6���a��p?.�~0�!�N�0��$5(�@�(�u"(�Y��H<�ђ���WO��9���A'�D�Ӵ°ԳJ�	���$�:�
	�%*��=���n���w��u]o�-�^y�����/��J� Ñ�s(a8�@�tX�N��<y���z+�$Ӆ��������H���� q?��W<°;.��/�GO���M�M��5���2���k��U��I�D�0��.���1@9SwaX��`���{d�B{!��l0,޿�����LX�m�Coܸ��@�DI,��a/����ώ@d��Y�H	�N��yI�� �z���Q1�D�Q�����uWΖ5��U�(
�<�=�c�����������b�9�ur����"@�k�Ϭ :!t�@(5���@��@������s E�z=�3���,;�ڇR�u�_��>K��R���<��U��s��;a�v����,���!�y���������s ��ܬ�}��8oO���<��y�\��9������s�3w��/�� �Sn���X>r<��c�X?���Ls�LL������%��\3�,l��J�A���{���a��L��p/ ,�ev��m��'�i�J����j�Mg}�	��G!H�ظD4U������[�p���qq�f\��#��j=|��}����O_�W�_Ǯ��Pڽ}�~�N�^���7����q�uX�d:;� '+����s G@��b����%K�n�������Q	��,�߁��g[ax�R��@>�|��{��\%�����o�įw�aGN�G׬�Vn!����s�R)���dJڑV׎�"��U�{z7v}��O�÷W����}��=��=���|we7�w��o��?\݅���Ə�v�{�sin_��]#��ڇ��=�o��wW��p��!p7Ϟ��w���	����Ň��Լ�dVVcf;S;�<Q�2R����G3�r<V������lǳϭþ�W����>nr�+���kp��e�Y�,La���(�Tbr�X̙<�N�S뱠�������z,S�#K0wx>fw��:=1��0k��@������>���8x	 ��`��D�3�\>�H(��y1�W��wc��ɎBB$���g�#����3.^�Y0��
�	���R�� |WW#�@�_}�jC��'����~m ,|W���8K:v��l��p aX�$$���H�1��C�h���L��'t�f�e�<��m^]�o�����L�:���G¹��q��I��z/V��B����� ���
s^��2`Fd��F�V�b	�	�"H�`87/�Ņȧ������B�v"a9��>���@x�QI��Օ�(.̃�dP0|�gXy��z����:��Y X�XF�+))��M�p��I�޽�o����f5�HA;;7S�O���/`���xr�c���@em)R2dBES=a�U��u+�q&�
���B+��+�F���}��$���������`X2<�`X��_���<����Lk�6s��2!�������	�˺Y:N��@}�P�a��
^_,���M{c>\�1{&<Y��F��h"��%}ؽ0�r��=�%�W��p�).�9|o�T:8+w������ĪJx��|�"_f{
�L������{UW�����y�9��<<�w���⸻����i--P(Z���;�a!��v��1��I����vr]���^:���#c�)PL����w̖�Fd�y��J8���s��އ�}�F��;߇�K����З��:��*�]��!p-Ǳ��m��r�#����-)۔�;�,Y�mg#�3�(k�R���Sp.��0B9��\m�)^�-�yuNN��hY/poږ�I�(�PNC�y[�t�1�۩�<7�Y�|e-�r%�NF^3+��T�dT�gR	��W�mh�d[y'��R����;��J�s��fY�:�H	���&+A�W�<����@'�	��ۄ~�
ku��W�&@v�{+�fI�A~]h\u�����T��R>�Ky�r���	��f,L���wU�v`��ʔ�u%�v�ut	*Bg���ٙ��"Fi��НߔY򟇎��H����"P,�$�(c��v+�O�P�c�� ��C�JG�p�!c�~l��J߅�m��|��Ik��5!�J�h��8^P����:�����q�o]	�I��!�����O�d�(#mv�Ǣ�G�����������G��`��%8�g-�ވ�?���:���=��]�����A� |��SV�ľ8�g9����v-�E���c�p��\?��mŎ�K���w0lh/�g$��P*2�ߠ�G�uI��t���i��&�H�0�>��͝�/V���3L�Onnz@�����%fX�X@��_<~<{���	յ�0z�G��Q�]h	A��@L�L�{ƕ�b�
0��9�d+�\A����pn��û���&!����u��T��m�/�����d���<�ޣ����2A���=�A@>����A��h����"h�����7n"��R����|�3����8�db���	�2�0�3k(�&bӁ8v����AJj/|�t��?��W��__|�i#��j��w?EhT.�3�3&���3�Y}�����B���/ƕa��r|>�����{#�P��_7����������N	x�>.��`L�����/
��'S�	�x䍃W�V���W���\�G`.��v�;��Y�J	O��v)8��>/K2Rh��=;��fy���y3����'�GDV��x�Xس�w"��g8���P̯°3b���&�T֬|mC�56ɕF�wRx�����ӓ��Ft~_�<c������PRZ��,�\����~3��jp��a|��ǈ�����-�|�K6�`
��&�ʺ��0��F��C��d������X.� g��"1>ɉq\���`4xq{_$�E"=5��wRS�wWg�:�"�&{�z���n.�j�鮅K�0�~F_�p�^��p��a^O=N�:��Wo���c�2u:2hЖ�Wb��Q8p� Ξ=����c����vɷس/��`A��k,]��>_r�/�_ᇍ;����`>7	Oq��J]�p*�NB�FY:n	�j�!�r��	ԬC�(B$�W<�rl	P#ظ����FB�L�^8v����
���|2fWßð�إ��5�0��~�$�L�}Ӑ��5V~�	Ȅ�[��Ip���|Ig%����n�sɷm# �/��H@ؚ�Ȗ��)�
�����SӘ]�l@5U�,t���(q{]J�$˛ߙȓ�\�:�:��� ���+r�rW�%�?\Y.�̛K�d��	뢶�x��g��Ã�� �w6�n�8�%�d�E��:�W��2/�(�F��h1
dDTN#��r��6�<~������5~ �nO�É�䭶�|ٽ�[R���fk��G!Nѽ8�NQb�h�e*m�(�Ǘ�g�-��e}f�c�q�h��r>;����k1D(+~{"1J��CCC�#9��:��O���y�Q���>��@x%�S��B�l��]�����t^)�H+�|��o؎F�L��L�0��1���es�q�X��s6�ʻ;Dy���>�*��-=�و��ɞ���94>g�3k2���L���X�M�[-��,m`��-��?"�T���'y���N��a%uAX��tؓO����C[��DTr<F��U+��٣�q��zz�*\&םܢ��&q����[�3����p��8C����kMZ��G~h��s��|r.߀���b������)ρW�?���pKc���z�64�%7�t�����U`�ߢt�sJ�߂���L/���aB����G	+ �'��_�mҶ���#��c�WjnbԌ�\1�UV<�����9q=G ���S0�ݙ8~z?{M��p��^ܿs-w��O(������޼t�Ε��}�ҭ�^���"�4W�'��<�_�g��p�<����n���52{Ν=�)Ӧ����T��O�_B!Bs�#�l��&#�h<�rG���X:��^�����2�Kd��øI�Ĺ��T��W�Ǝ�Ǳ��!�:�iUHH�EeY%�L�����ߩ�'�����B|:� _�/�WK�pR!L.��19�H7"��~ޮ�%�tu֡�c8:;���;A/z����Ϝ c�d��O�o�DM���;NU�݌ٰ	�%�.XIxr�����
��a�� |
f@Gx��\-,A���Z|�뤅0|s_��!fu�]�L����3��(b�tg�ʬK@OBL�ܞp& ��Ý0�I��,�°��sD9�X��� �И�ʂ eG8pae���U�b�%���7a�;���̓OL�rhHe#-� K{;[�bɢ��v�
,��s��T2Ҡ#�:;�#�@������t��ONIJ$�)�Vۅ�!:"!�@H�b"�ow­+�|������45MJ��9	�:/�|���Vϰ�Ix�y��U؄��3\�\���b_�QAsZj
>�p.^���������l2�s��r��_�Ͽ�c0z�x�?�clݶ~�r�1}�|���	h�g�2����x���ȹȽg#-Ɗx�;�p7��'�LV��1��JJ�<T�-�E���x	i�Hf�E�
<J�S<���z��{NDr�wU�����+'��⅒�֟�'��Nw��a��p�88�auH(�`��;�7�0�1^u�y�����/C��덀��p'K^_��ſ��a��!0,7d��Ar$��E�*g���H&|E�"�´��.&�;ϝ�(��.@/P�A�Hy�Mr�u
*9�c�"�8��S�K{�C�Q���s��;����"G�'p�F�t�u�G�ݒ��Ir@�p�*^o��6I~k�p9�7K�% Lv�u)P�fu��q'*ɽ�	Ǯ�,K��7�M�<�\��G�E]� �ߑ#��&�9�g�m��L;J�.#���zP2��J��%��������L��\���v�:gʅ�4�=W�\30Ԕ����ܓ(��E�[�]I[�>�W)ܗ��Ybyq�Y�ʠ�G�W���i[Gyp�A�,���^<�W�@>�����]<��t��xf�#����L��J��*��z_�
��\�4K�W�@����"*A�3=d���!�ǬG�it���?~Ap�7����q���w�o��;l���?����8�s��]�+����M�~t3�ی�㋜^���G7v7�7����8�mO�O�O|O^�S�W���q�����/�{n>Y0����
�k`8��a�/Y>X����F���e7�_d{qf��G`���7{&>_�=>Y��v�$t�%LB�DwG����}4)(�o�៟�_<Q0|�FFΘG��p�X�ULAT�h��DRa/��1O@��46�D���hn܎����=�n��mS�Ԟ?�+'����è�p5����s�q��~>�]�Bv�̑��|nU�YS^4�������uB�Mܭ;��O��_���(��DxL��"q�I�J�@t�H$�OEt�$��hx'T!,g>��G�7�.��ʵ{1f�<|��J��v�o�Ƶ{��v�N����J��*��1g���@̛Q����ө��E���pON�`J>a8�FD�[�����/�v�ƛ.x�C�)G�'k*t���aC�$B�h"�a���e����C���+*ߜqld�h0\Hc@`��Njj$�@��`�w�x}��g(y�	�`9����n�+�ە�v1I���m��^��saX�;t�D��	X�iG�Ty�;��'��G(����J��-�WD�������8$�tꄮ�ނ��%�(�υ��3�w�[k+��<�f�=Ĳ<%9�	q��$���S�}�����P�fe E�	DXP Ғ�M06¨�@h�/r�R���LHMD~^���DE�}M0�kb	��&�{{J<���aG8����م嶆e����{��`���0˘G{�8y����a�HHHGrr�ww#����g_Ef�.��xX����,R�ޕ!�տ��L4.#Lp>��-��!=��2��{0ð��� Ä>S@[�O�C�q;<��N� QEF�Ù!�؃ j���x� $���?��[H�ò�Q0�>^y��;� ����d�_�mS	�\�8T�S��R�)#`A��x��9U1��u)�7�j6��`� ��0�G��!k���?=�4u��Sq�*ƶ�T4�-]�9��h]E*W�s�\e�t��<�'CX˿��d�������(��T�o���&���Z���[�_��g�y�e���ȿ˥#�ēJ������ �*��E4p����<��ce�9��*X��\o�W�$9�v\��RY�P�{A,���m�j�$e,R!=&�	�C�,��T���\�PS�m�5�0������4D��t��?uM�g �(�{3I����x��n��,[ӻ�����˵T�,?�k��!�B�F�so��5K�Ƿ�9|��V$b�!�2��pӠ"2��hؼ��+LI�� ��*+pgy�8o#��ıݣah��H����O��N=���?��3g���8�g	����,��#kp�`|�`{��z\# _�.Q�Gw�Ƒݫpx�*ۻ'��q����������8u�[������-@���8vb->�r:�Jҡg����2(����&Bw��Ȃ���� A�����*�+����w��{�Uj�OM0\����'Cr���(���IH�|xz9��Şcq��m<xv��^�&�4�������(�6����x�X���j��v-Zn����;���	���Rz�t2�Ec�UT�=�c�v�a�ƥS�p��޺��ۗ���5<o������:�<��{M�زub����؄lD&�#����ƾ�$$�MCL�d���$�샧��5��'���{>������Qϛ����{�4���~	���Byy)fO��釹��yS2���<,��_O)%��	��rJa8�2��%i�Y����G �t��_]���W9ceX��Ξ
���Jf(��L�Aқ�Ӓbc%�EgV�~&�-�C�4�f� �x�ۼ�S�C��I�`X�j~��^a«�`v�2Wʙ����8��"'���,e�ŭ`����%��W`����`�ܟ0<�0<�0S@.R^I	+y�3L(�-S�a}\!�#��O�Px�`��CHp,�u����N�S�`�`ce�`��׈ )�c':AS�JH.त$v�#�B؍�'�z8�1���DBt!8YiI("�&Ą�����+���B�hb4bc���b�%�"�� ֋K��:zx{x)���G����`ggG��:wⲮ�ڹ,eh�o��m.��e7[8ٻ��۟�	+k7XY��GB��o�i'�P��b��>��I�#0�������	��j�`-х�N���	A�w0,al�%o�x���&Q���ᔆU���߂@��G��U8�YK
68���{b��[V# �\�UB@O�{%�W0,��lU��b���'{�Ép� �Rd`	���Ü	�m�;e�U�M�4ð��t�{�_0�@=�i�N`8B`��B�&䉡+�lL0��#,��1��0�.�<[�iH�e�:�@��\����
vy/̙T�4���d��RK��,f�|�a�̙)�J稗�sܚ�Q��x�xZ��ujn�������Z̒0�v�ʺn4D�q"�[,�\���E�q;QW���&sgB�����ԍz�����Ԟ�C;�2*��:�΅�1.[I�ղW��k�Lb�^N�:���;�$!^���Lei+���x����:�{[��N>�L��7�C'yG%�t*4��)a ���c{�*��'�$�G�5�R0<�Pi�"1�w ���`"�a� ��rd����N� ~	�����\��gĻ���Qc/.�\�����8��[�ܳ������qb�
ߵ��
�v����˱w��{lߴ?�������ƾ��q��� P�<��0�a�\��.��'����S+�g�|0*ҋ���HXI�5�F�D���"y ax\2 �d �ϙ���Ǘ_�=�v�a�>��N����3�A��;�~��&��a�t��	��0b�\�TEj������q�/����d��77��Y=�_B�c�ww7�q�����N�G�񢥖���[�������o2����(?~Hx���O�y#n���7P_]���p��Y��e<�w��}��_������x�|���b�� ,8��HN+Ept1l4�� �|&bJ� �p��c���\]+�?�Դb��`N��Isp��5��ժ�((����HM/Q0<c�`̛���?���Ϧ��6�/����1xotzg�!��g�pw�[��7����l�ջ�a8g&$�� �'��� �GJ`؍V�����j.l�\ـ{'D@�NeE@&�
���t�	�*lB<���b�� �e��N�I6K��m�W3�
�:��Jaʅ�.<�Yn
�5��L�Q�qlgM�ex_V�°��0�ĕ���a�7�S"4gax@�	áy���L��mO( �EU�����$U�_r/⋡�̄�4���}0y�T8��1�HI�ؑ�1j8��DV<6Vp'	���M�0,��ud���tW��bc�E�5�(oqDX(�zA�Ѵ��c�P������e�"1.:�;�����BBrfz2
�U�FP�?�����r^�	�>�F°�� �{����{{t����b�ߖ@�Cr�7�{�����ڞ��檃�_8���� G'=l������TxxE��=�^1�r���G<�{��!�� W��^ M��\�`�Y�བ�bdD6}j�^�B ��"{e!���g�`C,�b��C$B�F`��g&P+�X��N|�*�4��(�0�ӆ��ƒ �x��_��ے��x���0�����F��$�I�_IG�)m8�X=�%m�*Av �K�5N����ǰR�`X2X����7���p�퍀��peCm�X}�t\⵵fy�+�@X���2���0,�ģ&�D��s���8�_ 1L�V�m5��7�������	u�N$σ�I<�bt���$��"��B�I�u|�<��m�#�.��J�YZX�x.e[�tjS�Sd}1�l (#@ R��O�AjG��&(��X~sJ��m� J��*p}�Y��Fm�2#�������U���p,P-�#�I��v�B�vlQ�c��j;�~�s�"��H*<�RN��!PB�`�^���+��fIjC�0�1°a�J:��-%��&�MB@8���!6K~|
��C�U���NnU�R0L�wJ!HVֱo��J�c@(�89 4>��O��C+Pse;�_،�'�.ř�Kp��2߽���{W��э�|r��߃+gv�ҩ�z~��:���v�ġ�8�kvl^��/�Ƶ���GB��U�rj-����|�+�ұ�y���>O�>�=>�?م�� x�D�#6�qŰN�����0\2ߙ��֬��E�o�<n��`�nc3��(�O��W��U)��4�A7�v��Z��H����#��{��	ƅ���'_�R]-�<l@㣫h||�O������2Z����ţz<#?k������a��~ba~��z��?q����I��-h�u7���څK��|���7�=���x��>#�_:s{�#�#*:aQ=��J<>w"zN',�U�6�e���˷���_p��>V�߇�������AX�k/A��.Gv�$�Bfv%�J{*��3���ܞ
��3�ax����y#��ިl��D��	zw't'�����%���Y�w/~̱c�-�&J'A�7>,�x�uY����+aX*v��|�p)�#+`L���+�������X0S����ÿYMg�5��!�;�IL0!�ru a3�Q�A�*"M%O�+�妀Xӫ0,���������\�;�:N�E@�0��a�a���pd��N8(8�"D<{��C�1���B�De�����4L��.>��S���@\T$�"#������b��MЕ�`��N�O���^�L=��)�!$4X�vvvDhX����G/�tH�/AX`8��i��H��H�&�����c#ø.��b����:�y{z 80�S	���	�^�a/� ��� /w/8;8+�ޥ;�v�.����۝`��B��-%�4��x�����r��  0
n����4~��π�?^~��ʆ�O*,��h��D�%��"��s*a�S��b8Jv��>E�证�M� V��%�y�ȑ��FM�5.�%nܚ����<��F'�D�\N�r�Rul^�=��I�b��*�x���d"�N�����ia
r^���.s��d���ð�^@�r��RG�.~��p����x�,Sh�~��fd�đp��!�x�'GA���S�$�|���9����0o'�ʫL��=S ,���C����}@֠�:`�,�1I�δ�	�̚ V��7���$��!j_��d�״������>(�p�jp�B!X'Ȁ�)�`�~_�%%#��,_@�:�cG�
��wGP���C1<�L��|��dJ�6͛����g��Tn#e~��z�^#�?4 ^��S����X��y��J<�2.^9�Y��(@�cI�'��dД�x߭#�Ԑ�n��Uv+a�T~[�#`+�l�#aW�B(�6k�+�`�K#Ǚ����5q�����K`�{�5Ĳ���>��O�M� ��t�������.�F�7玮��S�q��2�;���g�-ǹ+	��%bNZ�+��V�Q4�9KF��w/�n�ܭ�Q��r�<�n^"k]@ݕ��|� x;�ވ�[W`7����ը>�������_������q��'�xl1�X���Czv����fۛ��r>�>m0�l���＋EkW��o`?a�IS#Z����������'���	�G�S+!m�$����J�0k7m��_��^k�^�������4��Ӈ�q��1<k���-���p���������E���V�@�C�q+�m���-|@�Z���~�n�vmj�/���<��hm�ƣ�+x�z�N���6�`�ڵ�Hɂ�w�y�cz#4y8b
&#(g4b�'�3�s�lF�#�{Q�w��� %�?2{�ø�s���ql;|#'}����HJ)FQQ!ax>}o(>�U�/��i�X0��T��	e�xL.�������''q��&�pwW���7ܣ��4�o�|~����O�[�8��$�M0,����&K�aؚ�#�Q�M����(����Y�+��¯�a�B�S�i5����yg�<�S,�fp��*"�j"w�X�<n;�
 O����[��6����q^���lx��9���������a�?�� ��|���G*��=!G6��Nl��^�"_�wla��Eht�Y��.Ca� dd"44�vv
DBt4�A�ӛ��t����󅿿�[�xze�ؓ`�A�K�DT�c�ž*�ZJJ"R��}����x#��Ch�� ���@�o2Se�Ӆ0�GdhA8�e�GXp����e���Ф�T �%�)�,s'�:�:~�ѣ�,��@�����o�o�w��/�_����oo�G+�⣠7�P�茡
O��W ��r������!p2���7�p|?��ct/�9�̑�&0,��9���	� �$�K�OV��JKu-����xJ	�	� �*L�r���d[B�����w��NJ�
�����Kz5aYg����Q*f�2X �@�$��.�9z�����ֆ�|ÎaG��#�;���BN��	{r�8���*D��/�c��a�p*��l�d�ϰ-��l��@X��""ⵛ�*�J�&Lb�%���Zl�mO������e0��$ޖS�6���!�c�gW���Iಠ�.R�z%�Y�y	UR@l��~J&�r���c�^�h�W�������,���$�u[�����6M2�8n�)t�`.����L "��cRr,���W$����fɱ_�`��uq�?�Q����vyo�P�-^�2-��1'�j��|�ԛ]�.��!�k�p���SG��Î�![�`�G�h��4�]�Oð�k�����l��p�!��O!��%�md6zx���J��Ʈ}q����bߵg|��GV�W���8�k)�X���6������f�1�_?��'	�gp��u��W�7��u��n^;�;5Wp�������?`�6���5����|'����sql�<���_�[�`��ሊ�@ aX�{��URX����́)����ŷ?��7�.��=;�0�*0L�`�����9��gãg�Ej�@�������S��?��Ο�Ͽ>FӃkx�z	��/��sx��Z�N���OO��~=j��k��ţV5�V1!��}!a�?��jj�E�遈7A��=�m�%�GM�)4޺�����|�r�8�n�/Oo�q�]L=.N$$W!��ot?D�K�	����X��0��4c���P�ܒ���k�
�"9�W�ŕ[MX�|��������a���G�{c�;�pJ��N���O�ćc�0wd�UD�D�/!���Tg�����&�9��"����J��x�s'(������	�A�--�+!�=R�-F�>�x�T��4	�f��pGia��� ����1�I�<�M�Ν�e����c�<�&��k!8��GΛ��Iڔ���Ec�w���N��Z��.�s��0��p`1�	�n��]	�ܮ�����`�FA��1=' �x���#$g|{�ʘ
��T�M".�q�����W7�''!73�P�;kX[ZD]T���8@��z=���Ky�	Þ0��!�����SRx��l����Q�!<����p��&��"&���sE�t��L&��r���଴d�e����^e��(W�$�C��`X���w؇ �GWXv�B緺P�	�o���7�o�� ��_�����o���%�Sv�.0�� �gF�����E$ 0"�iO̅wH���iTd��_�9������a�|w_����a�
K�B�'�I�$��x��9��B`�0l�wF�����6������G80o4B%�7�:�S�-��]�d(eANF�+�1:z��.��s�x�5/�S�(�&��Q������¥_��
�eCR�L���=Ϛ �Xq�P^k�Ġ�12����ü>��AX�Ad���0A���F=�U؄�C��vnb�3,��\OY��Q��ۼ�Ր�|�Ʈ@iH(�0�(��g'2�)f�D
���1V�B����	h�%ώ��&�׾�۩}$��&K~�Vm���,�
����jt>1�D<N�:,S�n:��n�����OY�r���;n�����_��$�9^'�&( U��d���C�?�����:���V��x�?��O�˃�ؙ����ZFT��C�t$�͡�O�dN	¶�G��$�p�?
��f6K��O`��Զ�Yz9ۅ�
S6<�#��6r ���$Cĳm�1��z?$KW��&���M8��k��b�8��ڄG��Ў%ط��z46Ó�Kh�{՗���ɝ�t� ꮟ����Yw����k�p��)� ��V_��W	Ţ˨�>�ڵ�Z��'����/q��G�~����ؾ�8qp-V.�����R0���$��o� ��i0�λX��0�͗���xF�k%��#��������ۋ�	ÿ(;�]�����#ѳ%�{a�ʥh���mo�~A��<!?z��'p��V\���W�����q�@{[�0~���.�S��Y�[xb���hi�����R�4���ڥʒyp��������ߞ5 ?�`���BPX"{�Y� m\�t0!<  ��IDAT�DT�X,�u�o?9��X���>H����"�$��E����V�ql����g�e`����ݑ�5��,ü�E�7��'��g�����p6�+A����ypc�j�7��7;_�����*o{��
����~5�S �E8�ɛ פ�
�Xq���ˠO� �sAؗ�i$��r}	�"�@p�t%=��T'9Mj�8B��a��K�L5�Ѧ�9�XB�!9g�6�����& �hs2�r�dj�<ÝSw����j���a�$/���p|X����(�m`O����K�A h��^&n��0	��R�e��g�R��f<ėNFɨ�P:z>R�f �@�9�1%���)-�gK~��w>ƪ���k�|��<|2oV�=֬X���.Ƨ�q�� ������K�5ð�S�w°�^���9R�D���I���ҧ�x�)/pld0b�B�H�99!Fe��rsBan�T��Nv��諅X�p�
���v6�Ix^�����:�:��֊d�pGhPJ�{b�ȑ�8a<&N�#�!22�j��q�&���?��ŋ�|�Z���X�n~ܽ߯߄�7n�̏�DpJ.�`�A�ɂ}4��R8q�)y�3�V�<ź�~`��0<D����V����aM���%�%����tː�"�|G�$n���� ��� 0���>S��I���>Y
�<g|�52�kL/�����p tv��l���<v�d��1NvIC���X$q����N��B*!�߇��(DNb�9!=�{h_��HH/t1X9���!kY,��vf�k��+���6�杕�Yb(�^6/�F�djU�A�����:mD=M��e�e�2q�C,`��/�����0��&K�J:$*i@��)�6A��۠X��s��W ؒ�H��r���sX6�{��Җ��1C&YPrlK���t4�:�s�B5^����}ݹ��_s��K�am�C�;,���D��k�`�N�`��A�K�B#�Ek������(G �L�)�!f�܁N�an���|_a���f�ǀX`�,��aXFϳ��e�H�n����Mc�5��p�6b����A�t~N�[��ǖ�ƙ��tt%j�n��]Kqd�RT�ق��ϓ�.�����<��k�q��8n\;�zᴚK��Jwo�@���5�q5A��W���q���n�����{�J���-�
G�Ǳ_������y�%ؿe1�8щ	��J�a�6���Y�dFH�`�߮]�`�a�ys#
�6>@�����/~�O?��+5�7�]��pha!�O���֡��E<�-�gy��t/�g��=8|����qz7n\>��[����r��.��֬�����$��C�^ ��+ }�N���ԞE��s���xp�u/]%����ЧO_��BS����0&�EH�h��.�/f/݂˭�b��38j6rKF"%{2�a��Y��n�{�)sB����;i��<~����KT�ļ�=�޸"|&C0O�����9�`J/�-�G��nV�u��[��x���#�o�x�=�F	\��C�9�����CGP�����,�Hia�[Z#��NFD�L^�΀!�,c���k* �����=6)��7�@*��"B�A�3B�!o*5��=��f�<ڹ�<�x��ܮ`�+�i�D�x��	؅���Es�=gN�]dX��î��<�&V�n�
�n�ᰜ��K��ׅF�!�0�;�i��b�u���H�5C>D\�Ij{Ϩ2Z�4��©��}
�޴7o7C���؁�}���Ϋ �g���r���k�!59��16�M�����I�T`8*&J�<'��:�QB��WG;�	�������(�G��p����)����*n8�ǚ7w.fM���%��K0�:�Ib$������nNp�w�����2`6������z�u�x�<6mڀʪr8�8����~��;�`��}�y`�}�1�[��׭�����?�ź]{0z�{��Hj�xYc	�q=	Ä�����W0\�B$t|f�0<�0<V�%lDi�s�d�ђԿ�|ߥ����2�j�a��	�m0�Iu#�	���Or�! {$B����Ր�bK=�n��U���&g�ƸG ��z$q��4S��5y5nbW°s�H8Ƴ�
�7�E�O��
����>�7�y��J^Kt쥼;6a�U���<!�84�p�^��D��`���D6C�&��W Wd���XaM� ���W���(�f/pGu�ay^��_�6n_�@����j�����/ �m���x�s�dIYJ��b5�o[�����_�0��[����%��E�"`y;�#Sʐ���(�R��(}���`�߄�K ����rQm0L��f��0,��%�%�Y;~[ni�h�J
��*<�6e$� �o�#[*����_��q��@����˲�r�^�?��e�2���.�k�/FÚ��@�u�0����o��v���.��Ɔ����-��q��Z�k�V���:�;���~����a��ꏢ��q����8H>���QWs��8���W��h�]E=u� \}�
��:�ko�f�m�\�AS��ߺ�#�wa#�w��o����G�IY�ĮŸx`%�\����ĥ�1��|J?ؐa�h0<�w/Z��?�߈G�k�^�5�W)��� �YA���/~n�sz�����_:��6x�
������¹�{� ~{\�����ݓx�|�<��ߞ\ąkp��ܸ��oG� I@��ţhi��gOZ��`+����AX�H.�~�܄'���w����W0,��Z����)��݀��7o���#>wa�
~9CQ6�ɽQ8�]l<U�k~��7�r�Q,[s붟��ڻ������AV�`�x&B�����7{$fO��gs�ᣙU�pJ>��O���bΘ|6k �� T��.�'w��B'+wtsſwCW�Tر���c��� �*e�d��a�B�`��:��tq}@�80w<|��A�>��?�p��+m��p�<Ө�q� l�<y�홡-�L�d�nC��3E~��r�q<����'P<��̏��A�>�����q[�C$��P��&��v"�(��	�1pN�F� ��F4�@ņڍ��\/{wWL������h�aa�OB_��j�a;���"$k$�y�G�����7W�GdO�� ��Zq��	�]���]��ۍX�|9�Y���u~��Ho�Ņs���%�����F_�|m���������c㐞����J&��0$�ŪtΎjp����$�Ʉa�L'��>^��Q���v	�Ѩ(-E~���?��	�u_���z�&aT^awO8;H�aw8ۻ�x2p�?���-x�|�o�Ė-�1s�4$'������Ƭ�������w� ��t���O�|q�^X�};��=�Ē^�X�+��`X<��
���.�*VkDj#Vɀ �|��N�	�7+�G,R�K#�8R*� $�e����t/���?O�p���e�5��@j�e,�'-�pw°��!i����=>�]�;qfc�ΆW�$����X�7��Up�����^����>,C_j?X��}� B`�ٸ�`�F^�y�0�
�M ���f���,��æ�*��$�G�,�S�+2�<�<��!�o�̿����T(GI��%��έBI$�I��u���F���O�p��(�ym�V��+R�	�m ���W��'zwy��c�{�}UKJ?��K��۔%�e��AlKF��+l�aKB��@�d�h�a����aX@�eּ�� 8�e��N���r�'��1-L�V��ܦM�[�`I'�#$��}�8�>�8v��>��;���I��cԨ��|�(nǑ=��́ŸtD�XN ^��`��/p��f��>�kw���]�^�W��gP' \K�%ߨV0\G]�v	W�/���+�����;�u���kjQ�Wn�á�۰����"$������m_��ޥ�vzޙ7�I9��.�kƠv���A,#��ax�6���	���*A��A�!����56-�Y`����u?k.
�E�!���Ū�_�����+h�ً�w��y�I�����<����B��8u�G\:w�p{��x�r�[	�f���2�0/�U�ċn�������q�n5u��4nU�����x���o\���T��&">�?a���&"�r
b���q�Ī�Xw��=ꚁ�������ٲH/ ��T��#$4��"0<�0<�N�/>�O�鏏g��'��I�����]�/������]a��M�;Z����X:���/����88e�*�OX�UI�	�Yɼ�Ћg� g���)(W�+9G�v)Q�ۆ�z������Jva���/Շ�NoX�U�"�BS��VI ��ܚ��p��6��Բ�j�o��^l|D�7ɚ kBȐ�Z<�ˣ��5�eV��eZK��2��[?nK��U�^�ʯ�	V��X�:�!r	)�{7��gt��q�T'���Q��ApV0\��W��g؎��qWBP@�0x��C}.����e�9��A�J��U�O��z,Y�����ҥ�U8��~�W��V�MT_�ƾ=���W�"%)n�0H�>F��&/�<�t�Brj223���p����t��Q��x�=���vwFDH ғ	��	��@��R���� �!1>�j�e�1�y�;�VS0���/��G���nΞ��q�����K���i�ߠ��J��?�[��%E�HDD�!$"���	�&�7bǁ=(��eT���(���iS�݆M�j�z�V�}N�;'��"8Ǖ����cv3��i��HC�2X��e*�!����!��Q��.�}$[E2؀!ن�D�b�mJ8��E��)# �	��|'\�z�a^�i����=I�G`�%��U`)W��ɓ�W��� L �H פ��!,w/t���'~/]=2a�S =g���p�׸a<f9���Y��V¹1�\���`X@8�p*�K����p
�J��aɵ�zqY���X6�����S�⎞_5�I�	tE2Ou��R�bSY�۠NA�I��<�"�2�5	 �$5�%��k@l�a�,wW����
�0�Sv��aԳMïz{��]��d��A�OYG�6�j{M��b�)�N����q$s��u��_� ���c��,y�%�Z'��KR�ɶr�*��K��ҵ
��
��/o�d�߽�эߵ]\?8�W0l�4�i�a�*!#	����1�XX,��f��9�@�]�0L��ז�I'6;���6���̿��G�xs��c�c�=n�b�_b���نl�F��sry4�`���LغE��=�� ��~�
E=�g��l����ȶ�pl�\<�Gw|�����WwW/�F�Ճ�Uw���Y�ZO����)A��U��U��U�\�F-��o5��qݸހ��jQ�6�j��\s��֝Þ�k���R���Y��*���sqt�Ǩ9��\��
���;{ ���F�@8�BP�@Ë�`��	���6����HtM��>.3�#�)K6�4 p��+����`Y�a�2ax�����5 9�PX���n������p�k��i��t�8~i9I`-vm��Omı}�p���6�ᗟ�\O����ݧ��	�?zB=V�~$@~�J�my�y�%~�7�t�#?l��GM79]��0���
���9��/�p��!�����_8"3��R��a���7*&�H�Đ����{�ט��&�]��?^���s�����Q��L�r�G|L�N�ys�c��rLY��g�{��0sT9���'�S��݉�PU���~	?A�!�s�D[w8{���^��M*Dl�@��1<�	����˛ ���l����6�P��Bsf�Ć��@`�JZR{��T�ʊІ�tα����T>��a�")�D��_$=���(��M�%�	d�+�e9!��Aշ�bK�PbE�c(h�ҒoZ��o�d�FT���qz�$�Jʫ�F%D:�HJ'6n,��A��h��B��������Rx�Tr��ľ�`Z��1��@\�u��3���H���%��"��U��%����@P��H��_����c��m����1vS����5�V�V�-��� ���'���'������>���\n�� ����Blfz:����q"�|�z�%NM�Cvz��Y�[vsqB\t���� O���OB��|�`J�S��}�J:#��Õ,rw������>��w<�.+�T_�Ɖ�'��{s	�����ĩS�s�^,_�|>�-º�[q��lٻ�'N��4
��p:y�	�a�p���Փ�G��+̩�
K�x���&{$�U��4�2ܪg� �t<�{GC�	���!��!pK �R΄U7B�%�*�	G��E�#�cCIV l�a;���������^	B��W���Z��U�4�Q�`9�L�fcdC�іF�]xoM|�����_�-J8-'l��} M�b%��*�E�k�`�moIȖ�Țߖ�Á崧qۖ��YĒK�:� Fش$�ZI��R�o^D�Y��֞��^�.(�6��xY</�A;��vq9�C%O� +�`�)f���p���X�j�A֔d����g�`�S-T�u�Y&�kF�'U�s��4�͒᫭�s	�4`���٬�D����n�k��w�~f�os\�&)�Y �Kb����$��K���S��5�֤���� P�ڽxU
>eJi��������Ӥ���6A T���"��V�yJ�w�ݎ2{�;���A���m�l�囍�_�C�rJ�?2���kfY�[�KZ7��m�ڞ��o�/!4D�X����Ú�C�Xئt%�`)�U�J��EM��aX5��_UEx�"�l	�Ή���o�1}a���$�~��~��=�c��ᰎeY����=a�EW��% ����Y69�5e˲��d]� ��Xx���%6�.�JKĎ�Qwi�]�kg7���
��.�Gw}�����d�8��Olǝ���S+"���h�'׉��5�L��TG5���f}=�m@]���N�kQS5盗�'p��v������)m]��?~��;��qj��1r\�C`���ްI��]v��uҁnv����n*�>c�f �?&k��f/�k<��6�I[����_��1v���F~Y?<����Rw�7�r����������س�3\<��w.å�{������Ϟ|?���OL�`���a��.B�0X�FP���	��n�6Z�h�{��'�����'���u�6\��������b�V�?{bz�D|�Y�,�����0��D@�Dj��%6�J��pM���H(�������Bzr&���>���_��￙���Će�뇯�k��Bkm��o��'�`pU��p�����=�CB��C�n����]�42:��H��A���W4��I�N��h*|rFi�"V�N���S�N�pc�J	0:��t`�����|�cܢ��$ϫ�x��"�P6�&9�"'6�jt;n'��\� ���� ;����0�AًX���##ƙ�#��$G���y@Á�*�WS�-e��O�٪�1��ȍ���2<�z�;�/���4�\_x��%Fh�3�y�,{X9!�?�sƪ�s.Q}4V\�	�"�{D��;�B�q�u��;*�q���GlR:���Ϊ�*�X�[6o���1��[[�8�<�
Bu�
�}�>>��@,�z	���A���P0+#��*�Db��TALD(Ғ����r�P�F��f�NF����Bll,��F�S�XG&�����d�	���)�����4Dɼ�i�f`��8�<���"���w˿GIY�r�g�L�6��@i���5h(�L����
g����\������^��Y����\8�Yz��w���ST+=B���G`�#����j��A�����=��u8�����I�&�ȿ��� :�T�JaIYE��m6�����Fg6�]�m7���O&AC��o� �@IpQb#*4�+S�a<'�&G�oF ���+�[�x�=]|$�X<�"	�(�pD��/@go���vl�)�r����a���p�s��!?6�FB �J��?�WH�]:��AXBD���G�c�,Z2L�DȔ�l��/@��6��%0���w���&.k�'��dXm9�@�x��-;�p8������Ț�� 6A�L;��,��i�������+}h l�a�����w-F��vde��c+9�V��s�`D�=k��v�5�0օ��s�(yo���{j����$�l#)	ס��ԁ�"��!ר�����ȽP�,��Ѳ�z��o�&�7���R���"(aNs�r@P�<�>f�#C�Bm������ �p��m ��)�(*��I��RN)��#O���{)��E%l���r��0ܙ�J7~�V�}�� 86�,��1/��&B���`X�����<�[Q6I��c	�d�Bp$f��ۮ�tt�'ӨM�e@6�_��6|7�#����6b�8��0���r^K�r�;�p[X�+0l��J��}���@t��s����@8;�`@U>��^��?��5�|�:�g�/��}ߐ�>Ŧ���a-���p����'��!��@�@�p\W+�@�A;�1��j�m]-����� `\���5rV5u�.�ҥC8�w5��0\�����oP}`����FLb<<����˺9��2�/�J�a�;3���Մ�رy#Zn6�x~	�̈́���Lu�6��?�/�#������~��Rۀ���Evi/�����Sq������ǃ:®������\:��}�3�Wa϶Ÿv� �}O�4��Ӈx��	�=}JX�� �����7�ac��2��$��q�(�����hytgL�wPBS
��>iC]9�}f!�r&�zN# ��O�h��Bp�H���B./�ߜ�H����?[�U��c�7˱j�w8ut7j�Ƶ|�j���-���Rl_�-6~�k�@X� ��F��N6�*���K ����]z���}�6b��? ��?�{�X0>�=g��d:|��1Y���C�"hx=9�`$<��(\���Y���X�d%i�Vٰt�+؎r��]x,��r�Α�VN���	����QILW ۞��H5�� �K/v\N
���w����p�5i��[l/x%�cX��
����K��Ć�3���#m�ܓQ�`�x�Yv���l@���Bx��<����I�ζ�p�"�z�K�n������/�K+1l�H��F��ҖP���p�����,�Ü��}LSo/ox�{������A�pwuQ����P$r�UG9�$'jD�����@`�i�Jǻ�sNN;99)�6�0����|i�y���ݺڠs't�܃0o� $$$ /?�����{GWXXۣe�y�?A����������a����܍�%�#0	�$°x�r�<�='�;e�z~S*)���= L���/^�R���9�{�T�k+�Y:�%�&l2�m����!�F��#u a�'���Q�ؼ2�1�
�	���[5L�@����A���'(ۊ��k�	Ȅ�@Q9���&���@��on߱���o��)��ȍ����W��e��XT�h@��!�TȄ}�G�=¸��E�J�0,�{)�.��06�\&��u�
��0���28�ʔ�^S��πa�v�^�V�f�!ߩ������`�Z@�j��Kmۦ?�a�9*-�T�I�
�V��HX�6d�I&��%<�J��/KI��Z���1$��x���Y������v�y>O	�ɿ���3uq;�>
^y>52��|�Xh���#�ă*�Xu�����Tܮ	��P��e[�W�D�����!ݍ��\����o$���t^�Cb�;�*u���I+�l#�+��G ݆ﾞ�+��]���x���F��K���xC����x����w�&a�8��+�U-^�j�z&�r��C�A��M Y���`�yB�s�`�k,#�)��L����7V�85���0�`������k	A� K�E�(t��ҺY�<����ᢵ�
��\f��v�f��ᰊ�.�|G�y�@���3yj�nG��-
����~����qh�|lZ��lY��s[�*{�*�	µ���UJ:R�Xb����{��� �y.�E�Y_����A�6���� u�e46^Ǎ�'p��z���5ax!a�+\P0���G�q�b���'!��Ep�c[����^���n�Úg���K|�ð���* ��y~�!LB`��_�`x�;�#��B���w�Cc�9��woBs�n<��ϛ��p����%N�_����F5!�E3و��[���3<{�� ����g&~����T0��x����7�sO↏�x�\FsK����C�����4�Qlo	LAE�	�I،����^� ��l������(��@��{�@����'j��7�ڶ�}���؄#�7b�֥8�{~��c,�h
~8���e>ê�_`��~���!w�Ą�`��fg�;�b���y���3WPP5���e��w�dx̀�P�ϦUUE0��;+�T���)�d�3��>L�-\�����;��?,/[(��H��)��& �J�4�(7��-��:�e�"��o�^/ɓ��xPG��%SG��d�Kln�_]�+C�x����*��
{�
��g���"Y��J%��@%q�ne=���	��4�D��;8v.��stF�= �����\�d�#�0���A�R���me����S�.�%�A��r[�7�<�������Aj�9��ޞ�'������Um�p±뜛����R�~~~���P���z�-��$4��AHp$�7?�۹����6����������������ܵ+�|�3����=,�`��['wG�!*1�>�T0��8�O`,�!I�􋇫1.pf�.��~�#�>�CӠ�wAb4��J�@ #P9������wC����d�pO���ܟϾBA���K��r6�9��\B2���Jx���e�x�2`A�	��Ө!�i^BsfJ���(���� �@' (8&�Z����l��~��L�]k�JX	��T� �|_A^���݂P��'oy��.l	;��<�C`Ox��{	��9:���r��"��K@�`b#�&0��j�n:5 ��F�V�}xl�y�"xNAӑP,S�v���H�t7��W����U�>�y��LB��&��gb-�]�7���v�xє^�m0lbs�5�	&���~V}P#�z�ʡ�"���9��-Ϙe�{hé�y����Y�n�Wԃ����R��]V�c�p�#�SL�F����&���,��]�^`��:���C"D�55Kۆ�:���`4� �.Y�U ��h�=��c���||�|'nc�xz��<æm����v�Uy��$�>4t��m��Bǁm��򮇲m��Q��W*�➄s���~I��ܒ��4�ᓃ���e���!j�9����!��f �������k^X3�sk�eⱵ����4�NȆ�2��p��|&"3���H����H�gx:�,�o������g&fa�e����G�<f6A�	��g:��d��Q�����:���S`�&�v����wp��Aܭ�A��O���=_����Z7k�����W��ŝ���wj��kq� ,�UL�U�e��fM�J�&@|�S�\���l0Mվ�W8���M5��9��G6���%8�y!�o]�������x�v������Wt\��^����]X�!����Mk��ۯ	Û�0��.���}�p����u^��_�����Ͽ d4T��ϝ�̢2��ƻ�>������˄�h�مG����=��8�[���3ؾ�����K�a���f<~�Ϟ��>�`� �`��3�)a�1/��m0Lݿ�G��55�	��n�k	��h�K�K�Nt�G��t�-�<�=|����	�AP\.S{�;u0"*f"�b:��#�x
B{NEp�))��q,�&�(CL�s\_��4�:t��'�9~�,X�e�.��U��o�J;��7}��_��o��>��|�1��|F郴�X�@�p#�x�����4�X������C�a���R	C�X�I�CҐqj����f�A`�D���2��#�MFx�t���i�z�'!���'�����2���/����+!&E�M߼q�j��s����:J����l>x}�(%ʘ5Z��O�é�w<�H�1R�#�{e��g�%����6ɇpe�l�XQ�qZg'��!�a�-e;-LB�a�;}A��0^� �Q�k�|Ux�x�"J�]��=*��`g��o��!���CbR2����X������FC !311	\���x��e�7�H��%�RF��
���;�N�%��u��W�E$�7,$H)��O�
���W�r����"�$	�vuu5�G��<o�6R�@��6�}�����n�w��6N���A�n=е[wt�ރl;{�Jn�h$�f!>%�Q�0E��w}0<�!��E�7$�a�0�f�+$G����C�0D�O���2A�����I<z���u�qB\)!� &��14xbK�\�f�;�0�G��(*�wJ9U�I��|�4>��,��|�y4���,GL\#�4q_�06bA��X�%r٠��BW���AH �0�`�D@q	/�~�H�A��K�3	"�fQ� 30�ЙO�[���;���ԉ�e��B�l)�(��e	;�!hfQ\��Y�ʱ��D�u������u��Gv徨�l�n$ũklOx&��/n�N�e	�r1�5�XɅ�w& ;��ކ�*�2�h	�"l���/��ͥ�(ÜW�J\3���r^�*�%���	�L'ׅ�ҕ�Iȕ"�+aZ?n퐎~քb�{��6C����S���
�e�[���$�`� ��8�"FWA]<42��([����q�fy,x_��Y�,���V��6�����p
��Cbk|��=�w�|6]h�t���-H X��	x����L��vj�h�#�:�o�������%��.\.�C�6�4�'� ��fTxsh��n�{/�ڕ�����$�&i�8�8,��9�6��
�;H��(y��r.}�P�Õ�,u�O�P�ӆ�����+MZ�+e �e��/!ژ�7i\v��C�0�$�$lGw	9 P�Aج�0l��R���e��a����I�d�^��}q�����O?t��F7{8x��	֋�^�&�>ZD��U<�8�P�8�0>��#Yb����V*-a�,�d�KJ�!U����ܘ�nv���P|��ܺ�g	�g�����_��^��5ؾ��[<��B��]�{�ܺ������&i�f5p��:Bp]��-Qm�&q�-��J7��xT�U�
�o�~�Uܸ|GvI&��8F>��k\ܳ׎nř#{0n�D�&��ڲ���6�'�wq�͝��?���%�`׏?�+��'�ه��I���0���@�I�Ŀ�%f�jM=f�� ��%�-��;�����.)�G~xk�6���{{q��Ī|Bˀ0��s\��_����x��1�
?{�g�m0�\�p+a���0����	��÷	�u�vn�+0|�O����<�]��l�c����*Ñ�3A��' �	�!�𲩈,'\r]H�{�2��>��3;^&�gO��{���{sf�ۯ>��aώس�{l۸[7|�-�W���������T�"*"��1ZOot�jA�����V����8t�����*�N��p�%o�T�>?C.��e-e��`��bBp�l�W�C�A�I����SH�,�`�QL����b	���g�o�Y�hL�d:�M������|J�(�����xE�?�������BP�lW�l�3Y���.NK�C��J"��5{�>�_R�����3�$Q!"[V�@<�� l ���a.$8���SP<�ať"��'*{�Azz:����,>���&!5%�E���э�)�L0,�I �������"O&��&�`7&��%T">.�ɉ�r9ٙH��EP�?�[����ሏ�GTTBBB��x+�@X�V�0����z8;����=�۠KgK�B�Jtz��
��F����-����c�S����P}�8���8��������!�`L��� 7�4�4�hxx$�.m����Lm$9itK�Ԉg�4N�2�CT�#��%TEd�zr$�:F��2 	�t���%��Vc�&�Ԟ�O+�1�^�9��ɆO|+�B%��be�!4�
y}S�х��*9/�B�+Pܗ�!8����/�7�3 ,{B2�p���M���J�WP�J�&Uq�zbO�&�r�J�'Wp�����������h�I��|h.A:� ���]@ff���`j�2���2�Q}�>�*ޏ��g1E4J�_�h)�N�	�ޱ%�Ǘ�:�+SA��ޗ�@޿>�z�IUܮ����Q�_)	�֛��
u_D�˶�~$s�6��=7/��}�����3v% �DKX�<[��$܃�l)k�u$�%ԅ?�AÆ -�Trڈ�Z���@w4a?��"��z�x��wxO_�n1bd����m(k^���y%u���	h�OC�䯦1Y��w��SG)�hQo���',8+`�o��O$�y�6�P��h�lͿS���J`�w��bdJ���J��;���d]�◥��uDY�1��$ܝ�A�PB?���&ɼ@�,u&�[�>YQ�ъ��:�lLBb�#�Kh�x��YFOIiHؕ�/�З��@5�K�dR]ซo:��ӈ���ԑ�%HJ���d�H��W �.��aXB!^Ä������}c�d�c8������;�C�������B�d "&���
M�KH:l�2hȰ��{̶�*a �7�0<� <�� �;��=b�N�W�l�򞕣����1�퍈�����	��w�̾�8l5NX���W�.Ŏ��ba����Pwj;������k��Z�6�+�5�K���z�6 V�^���/���p��U�\9���W`ߦ8�e��X�󻗢��\8�SgOGHF6W��t|zVa��3�j�z2�b�ں��6�g��dkU���Ј��m���>@���J����x|�*a�"{��;�zk7ax/a�V������b��/q��A����0��0��" ����a�,x+/���GMw�z�-��h!��[�-/l������W�����B���`x�	�'(�p0�8�h2
��?4|���+_���8�pߩ�u�2A�7��u C��ıc���/�|�|,��C�Y�%6�_�7��VSkq��)�>y[~܀��Z���ŪVXx$l�a�U���x���{��� <�A�+�R`�������$�����لN�i>�/���9�Jf��pk�!W�K��-�#��-�ᚹ�י~�L���ӉxN�p��^\�M_^'������8JyS���s'�;g2��'�$oY�}��)'��Tvt%�>{,+\I�F����Y��'��9	^v,�p6x���rG�7c0�R��7��\/6�~9��%��'�B8�\#������2�f� ,&�O�� ��ch��#4$
1щ*� �?���i|��0���K0,�ߠ o��.:*����8��֚���,���!--My�###� ��`X�� �?³�.^��sQ`lme�B%��ܹ+:QoS]�[���	���7�ߓ���q���u����.�F8{���'�~Q�
��[@
�3�@�É��+3����+��~l��@J�#JN�<d'��;D	H�/�����JX��q��y���TX�E��.�8E�;&�)yL�CPj>����J�Wd2�\g�ˠ��������Ba:1~�b3����#�Mi��˄N�E����s0A?4�љ�Z9W1+��e��ɘ���T��{x�r})�U���7���%�w�L �#�;��5,Q)б���L�7���
}B��m"�]����0�����R*8��o�*�ܐZ}�5Yb�d��<�#����D�+���^J"/0�F$����9��7��C�;Yxf�8^/�ڏ@�H� ��~5q���\�G͋�zC'�a	�)��~4�/c �Q��A0dn�]�`�$>|Y�)6�j� ���D#` �]�{����|f/��@��&�K�\�T�)�M�>�a���j�]� �K����ձ���1ט��q;�zI��<���6i �8�A�$ݥ;�J���G��g�Px��d�ȋۙ%�'�e�Wu\�G�H�Z��\S������\�LI���\���I2��eN����gh��v	B�^��Ar��m�(q9�N%�� ��><__�A2���}㹒d�d]�Prb�-�A�΁&!1�b Ȑ�"c�/#1�C��w:��͒k�-m8\3ǘ`x,S�� �e�n�a	e�����
G�8�Y��W�a���i�"\:�5���ԑm�f�{�ݯ����Yg9��:(��~�u�}a�8���Z�NCIG;��3��k���n��˂�!��H�O®�+Psf�X�Ҫ�9��N���]_`���i�l��n߂�W����+���bM�-�f�-�&%�`a���"<k n�0��ݻո�t7���T0|�0|�×o��3��sWD��0�C���x���,�ܺK�-�������=��D-���/����**ENY%f�Z��]��F��h�����Ɠ�]8'0�q>l]��k��C��V�P^a��3��0�D��t�{�B?�b��^Ô�WS��W`X��w-M���Q<���-BPt
��ٿ-L"�j6ax��f�LFH�$�M�_�;ɩ���"�0���%��	�[����	��`Ӻ�X��+|��L,�|.�^�!�	-��)���]�u��������^�5J�ʑ���@8&!�m�ދC�/�߈i��o�����^4ޅ���7����I0LG`��d}��A�ﲬ���rzn/���Q�D>�3�Y0͆�x6�=稩�/���j�.�T�s6���o��ۈd���G�<�q���ΟAc:��:�˕��7˨#��95�`ݗ��WHX�� w)c�ˊ:�/t����a�\��Y�-�
����(R0�#�*�=ѕ�6�Ͻb,��zq]�a�j��gD<R��������GkJb�z�"91a���������$AKo������N'���AD`�P	���%[�� NLJ@Ll4"�� �^ބf���ጌ奎��Q���]�_+i,��{R&��Mww����3!�]����7����[�KGA����Aw+X�9��.�`�D\r
��+0p�HdҐc����DZ�)��N�F�d�Ɇ�o�
��^���+�?��*��>�/zА��/T<�����R�!���W*O�Ep�$t6$�:8���
�����3?D���N͆[P��{P$�cSP>t4z���a����=f2*��j�8�3'LAρC�[ Q����V�b�hT���AC�u�4z��:F��k �1=�$����}���O0�����⁣1l��H+폰�B�Ġ�;�$���o$��)���y9��-F\a"�	�����C��%L�	��	�4B	���f­S0�;���/��m4\#�ad��ӛꃘ�<� j1|hD��2���$,��h1���H L�G��x�e�5(�匇�_�O*<C�y�S`o���W$�������/n���4\������s)��
-�7���,��Tr���9p�ϭ��6�+,�1�(�[���'�Q�c�1���~��^�g�C;�XA9|n�H��_"��8�#���&��! ��Z2��T�����!	.QE4�y��B������G	����@2�8�N�|7�(�3����4Z�6{�M��T��?���(ɍm-^�W$�]�ȿ/k�7��R��׊Ri���I�&5﫥l�m���=�M�?����6(v��	��� -��6&�9ƚ`�Җ��w_{®�tp%@;r^��T<��?ą`,�i��m}��]�9�P,���,X��[>�
�޺ܱ���TI�m�xX��W�+Wت����d����]� jV���p^stȀ�!�����"�W��c����uxt�4���,ƍ�;p��v�[�"XW�CX����`C���(�}��-�۔�I!�H��?ÖN~Hc[uh�:ԝہ��ǵs�p`���=�7��?��`x���݄�N����?��zBpa�AM5�TO�AX��K����w�\����p�� ��_�����V��΅8�g).\�j��G��ԊJ�G&.�`x���X�|)v��F���f�Tj�-��0L���~���[V��3������K5!��w��a;��Iމ�k�k�|l^9V-��C�	�����/�ӳ�x$�j��<@�l�ZM2I�`X@��\�\t;?V��&����@|���hm<�H n:�_iċ�b�����FVOV�>�V6q}�"��;b�$q�_�᠒	�/�c�l��L��<I���N��S`��M�J�~q��al�q�M��_|��]��V����ظ~��ف�~�W<��9Z?·�}�!#F ='q))ؼs'��9{�Fl��!�r6��G 3@̿쨥��-�!�� �l�j���2��@�t��i*�F��)�R`Ԭ�!�
���p�V�7�Y8��d/N�Q��U��˼�,O��Uyt��l&%p�]�x�}�e�)�Ή��*t)g#Ċ7�/��p���p��yh1\Y����%C�DK\$�~����������c���MA'},��������z�L�>��V_���Gh�܏����i@]�m\�\��.Q�l�TGH=�S�����:��<<<	��c/��:/O�tbsP0,����L�Դ$$�#� ɩI	���/��Ð�w$33S�=NJJRϰ��#K':�X��+�ac��rk+[8;�������_ �~#G��ʕ+�m�6��a6��	��۝ނ��V�[��[6὏>��K����q��	<~�W�j���1|��w���ZDЈa��B��e#U��Y��10��=�1�?�1ĥ�$K~i�[��z��u�S����C0z0w�F\m�w�]�ل�;������]��k�p<��~��#4?��w����{���/���3\o���M7�xɗѣ�<���ĝ��8�u���%��0�}��ʵ8q�5M����u<�ջ�X�mr����+�����,���p���ã�P��Ե�-X�}�͚gC0ްrDJAV��W�<P�OK����t��=� �wr�C'�h8���ڗ@G��E���3 �������U? �G{7��C0z�8^� 5�XW7��:^���l=t'��Åz^Ã�y�;�f�tu����j�aSfc�ޣ8r�����-�N�U�YF�p�FG��4
�J��7�y?�q��}��������oމ�S���ƈ��?�OX.�{����
��{�)�4n��Y����A�0tr���!ݸ��?�&x��y�H�Q�xayG$N�-��!o9x�\��=r
��;�-��Î���2�gBKG��x�~��䂰�t?�'��:9��3��n \�i���=�:{ �j��3<��}��D�@H���VA,G��Q�t�kS	���*�Օ���uj}P����RR�yJ�q����yA20�����m�(�M]��X^�+�)',��sQ�2M2߅�u�Aj��At���JC�[X1z� ��,i������[�$,�,	��ⷭ��.�%DA��GH�)a!2̺�IԪ|�F1��U=ޅS鼧B!���:�d�u���3}|���-k��aI�f�:VńZ�2��a���*A�#ڽ��@T�8XH�B�pا�P�����`���H���� \;�����������8�o����9��،o?c�m�` 3a���8$���Q������c֟���g����Uz��Q���1��DD��2t���;k����T��q5���士p��:�M��ޅ�rl)�m�����rIx�&4WË�7��*����@l�6y�o^��[ոu�2!�o���C�Cy?�l[�3����8�-��?��~������BW�nU��{ ��3Kׯ��5+�k�.ܻsG�v�^�75���<$?R�P�|Ϳ�'�Dwп�?�� ��>�E��*���q�q��n<����4�n��������n<kڃ�6��I�߼�5�>���[�J�o�P�) V���UA�������&ni����p��p�U�y�*�Dk�Y^����:zt�1�/T0�;
��3���l�� �pa8�tb��N�[�`$�7�>��l�ܸ	�	������˖����ŒE�v�2̝3�?�kV���y������_�ͻ��æ����(,+C,Ag��_~�a60�G�D`Z?�W̆K��5��	n��?v�2'�+kAxt
��)B���B�^�ao���w�,x��j� ����!�M��H^��xw�,븭�|�W�~��S��ĆBq�$t'w���yd�R� ��0�=BU����%���C�()�Ò� 0�+&�#�`ax ���9�Cf|���Zp�w���x�"�=iť�'�s�f�\#H�n���x~$df�)�pdD�� 5Ϭ��Tg�QAi`���,!��� �����		q���FXD(�`�7"6!a���������!�HHLDZz:�	��*dB�%����@X��%�����������zt��������`֬9�v�QH��������p�<�}��n�.���<l��#Ѱ����e��c�7��o1m���`�nي�	���(������)�
n�#	�����w�ƌg�hH�|q�D�4�l4)�RĒJI��I��>��Y8��<q�h��Y���O����l����CrVv<����j�#��{�?<��W���/�c���;7���	���Bzz8v��LPn&0�����a���x�p���q�M���[���yu��<�s�؅+H+���l�s-\q��s� ��P�׫�O�텚�9y&z������/����)����|#߫[�~��K8�=X����}lzx�oV.p7c��yl��Hݺ�1&��ƀ�>�.�u���?���ڟ��y����w}�O��~��o7�ߨ��;r,���4>~�$��l/׸��Y�a�c�\|�in��6p������p��3���|��G�6�:� �N�oT	���Y���b0m��T݌U�#�ߜ�>na���V.��J
�6�Li0�w��3���?6��c�;�y8y冺�M4Z�`�����}�E+�#29�����DRN��co���N^f�K�u��c����F�����ع[8q�.
�N�_�UB�P��� B%0l�d�6��`�ei�*0�U1��$��N�<�M ~��[��r�&��[�������8���r�0l�H'@,�:J��,p.���̱�JTI���PDk�ߒa��܃�O2H�l��c���;,�o�d�To��9�@�Ct��U`�:Y�2��_!��1pI��#�`�GfeT�Q0����ƙ�X`Xe5%4k0LM��a��`�:R�p�C=܂�����Ҽ�8-0��v|M������.G��xiv��q!:���������br/8���a؇@�A#��q	زv	�]?�`��ɵ`�;��>��\>���:D>p�� ج����z4��`XS-�{�y���F����?���8���ۿ�@�
���J��)����A.��>1��9�~�z�Z�:H�kQ�߻ۈ�F�W�U�������s��
����F`%��óg����a<�{O���-G����zk��Ū%a����Ys??e��3����?�@X�?�E����C0�Jni�Ga�~�y<�p�I4�>�G-���i���G�������2xG+��0	��p`�tB����)(��0�.0<����CV��w�AZRܝ\1e�$��~%��4 )��tsBJR&��m�6�A��f->y�{va��5x� ������0|�F�APZ�m�	�����ߢ�,�,x���&B'"�s&�h��+�B��@�IU�a�U��&3 ����#0�%�.�$�+�	�Żhދ�rl"{�.�7<�{N�oaX5���J���o.a8�0L @�����1p��R
�	��a�`�\4l2v���K����a���vl�Dㆠq�� �D~�֖gX��G;,��#lRB��`��0�}@ �\�!P,���o��!��b#@���`�&�"":A�A�owO�"4<A�j�a��
Þ��*Ä@���H�4�<�S�g�~���8{�,� o߾�˗/c˖1v��QO�����v��7�?v�c�~`�#B`�l���|�C�"��u�s�4��� �9pN�o��Q���p'�r'�G�.a z�W�Y
DH�z�
���M��k�I}`��n>	�����a硳4���'?������-���',l��W���7�n�Sl�)�O�FՐ�ر�������m̝5	��64F���҅��Ӏ�ׯ(�E��񘿚�k�s�>x��7n��q�Q�o���뷠��!Պw?��|�9�޼��}��;��������~X�z��V��8[]��GN���{���]�%}�ϐQ���EX�m��m��ǿ��-�K���;�	p2���; �y��g���iɳ9j����� ,Z��<ׅ�O�����n�n��/�0�q�f���/	���aϹe�a<x���k���'_-��}�Y�����v�ň�ӱ`�
��w�=��_b��1��.p��oB�~���d���g�
L��G�Nz5�@���O�9V�q��{�]:ЅJ*3I��k�dia�)+�dA���2p��ouQ(<�\P���!�o=O�ƩKl0I�g��c�������)����A��4g8}�Y����.F����׃6x81@���i0��/�pW�O�x�n�FM�E����������#x�p��A��K�\�ʣ<Ú̞�v�qXS°�_'m;_��%������<&�w�6Ȇt�sO�b�e�ub]2Y��3,�d��ps���dQ]�p��#�22s����Bw���Nq�a�?�a�	�G����Q	��MG�U�t�4J���?�P���ƙ�/y�O�ZL��Ԝ�G��@Jl0F�1�����ǲ��!��`X<���K/9��)��L#�]yp�)1�a�X��s4^;�`�≎0L��%axlX�s{W���}x|W:�ՑG�$����&���6�u��fnb��͛�`3�o�$߼Hv���,NY��������xx.\�+G7��m�t��H()�'�mC� x��0֟�>����~ĺ-�q��	<##>~�Mm0L.$������&����6�V����3��7 ��ᬲ�X�v!n5����W�|�(�4��q����/-'p���ع�s�Z:��g��E�:<�B=Tq �	�O	��O���c��0AX�����wϙ`����<��c7������Y}Pb�+�[�H��j�ʦ#@R�I繞�͞�]2���	��;��$T�Ǻ=g��������_o7/L�4G����k0u�x�˿��л����ܹ��d�7X�b�؋m�v�an.Y�ܞ=��@�b��"9�G�Q�L����Sa�J�Ț��> �j�aM����;��uXS�
E �f�fd@;�-��e�؎ � X�|_'ɦm;���V��W`���	¶ô�CK&3�g��a��
�Ɯ!��r�hQ��~��vY�]�8�x,�i%��K��}ǰ��	lܶK�[��>�?�Y��뵨�р�o�0���*OQ!���{D=�����:oO�L�
K�`_#��p���Q.<2������G@��!�	׾>��������S�����@��Ct�&!iwwwXYY�y�C�O8;;+��X$��aÆa�޽�s��OK���V��-,,Bxx�ʠ�TN��W���-[0b��pY2UXR����x8N���^�	��J��·Kr��Ë�K�x8���G�8o"�X��'����$=�����V���&Y�{�+�����
M!����{����/xBc���i<�����v����<<��b�Jtw4�ʕ�2,	Sg}��v�=��o�Fr|4�S���M�������_���B,�q��-��v�&΄�O �X;���#&L#p]��O����!|?���;�x��-�����I��ܰ}/�W���W��r����!�}��_B�?����~�JO��!ޡI�	�Eqy�ߴͬ�$^�x��OBw[gxD�M{p�_��,A4��p�|=���/�YߐD�|���}���na��˵�q�)��MH�.D{7$d���q]c�]���.~���'Σg��p��o#�1h��?~MO~�����Y	��L8�&����*�g���Y���?B�Ϸl���w'��´��N�VU���/tɰ@���K�K'��1��L�h>��j��;�0��%<f)Bb
0�E�z��|�mۍ���c�ϡ�~!����GNW#%�V��)���w�v.�p��l�N^nDQ��x�)��l�aIh��Ԋ�k%�@;H�k�OM2*bw���S�p�GY�E�J`�Ed,����5�U�n�%��zL��+�؅0�9�Pu �*�! K����T��nj�Z.eі�y�����B�O�F����eTwB�x���2�x�e;JR�u��o6��աVr���f}<@�-�T�l3�]h {���1]�;�Y�����< V�3lG��Kk	� �J�+	�h�a��%\B֛���g�2ul�&�xc`?�����}p"��$�D���-h����.������5jz��:4\ڋ]�").��!Nd�����.��>�0lc���%q,��u,�C�H��a���|�D����A!�v�{�S�W��Q�$�%�[H8^����0��k>����QsB\%��ð���Aȴ�o�ð�F@�k���=�f�E~�Z�������5ط�+�#^:���,����q��&|��\$����`��`8��L���߱�m��3g�\�Xo77���.>�?�y!0������rͭ��p�B�b ����7�j�1���7���]R������t�8������EX���X��}l^��.���G����c�L~�?����̄a����#��V��ĩW`��G��G�wU�ĭ�3�37�&�1����MB�"���AH|1³!�bbz�AD��ABy�	�*�X)��l*����0|Vy���ُ̔8�9a��q�r��\��M?�Ŗ��r�,��̙=}�>��1�[�[wl���\����s���``���e�~������w�;�O���Y�Ι���p˚B�$N8s�a�6KGh��a�X��egP~������+@�*����<���㶢W�e�����a7���4�0�?�0\EfC)0�[��!L0lC�u���![`x(��*	åp����c���*�!������'�9�&c�G����W`��OPH �<}6.\��}�>Z1�o5���+X�l23r	�F����X]-4B↽���o��
7�<�F%��� ��u�3�cЩP� �-A����h�ZdL�Z�Ix�&d���wE���2��2
� rPP��:ѧO(���T'�����`�!�?�oT�#V��?@������*�xȐ�6m�=�e߯����1��ػ��_�������w>ƞ�g�m�)B�7J(��_:��s��/^#Uo3n���qy�Ad��%v [�K�D)f8M=���)�����*:swZ������ޤ�~���������'>[��@�>Z�<R���ѩ�4���� �7���W���w�QW�%��p�'$��ex_�'���k1l�LD�!�I�FrN��S;w�0��,\�KV(>s���T��UT����eAs���P{�E�֍��x��/����f�m��b�тŨo~���߃Oh�cҐ߳
��,C�t$y�:�����b�qp x�G'c��ڃ_0������AP]ߪ���n����E}p��\mh��'����庩<�Ɛ(���"��?�T74���&�ۺ��"�?î�'Q�w0����4#���U�)�<]}Ye��O��1
�X�tjo5)�������H/7�����_j_x%T��߬;�K���T?�Ӑr'�%��;�t!yH+�U������Q�{8\�p�CFa_���
�8{��F��W���˗�r]�򔟫n��y���*�9�}��?���k-�N��{(8Ni�!-#{:F��9Z ��s���JYV	;��/�.����m�8�&�]��`��sk�U����qy��#���d��:�dk^����I��Lg^.��L��T/m�4hŲG�|�TsJ�M4�8�n4*e�$��x&�w>��� ؅�+u��F'C����ߦξyJ](��le:�C|?8&�����~��H�u����:{���m�#����P@�s�('�9���$c6&�s�$�Q 8�s��� ���z}{�u��Uc�9r��ߚ5jR,��%:2*X�W�WD�J59�DdX!5�"�!���A�4��B�G!��/�_�?�[�28e �>Ĵ~�t�?��;�p���;�-�\�k�����{��6xz���'�r?�4�7��,�E�'��)��*�z�1��3���	��|������b��}7q���s \ƻbvs�]�Q}���͸zf3.��N��ş�����M�px�J�8�=�SX�Rl�Js�'xB�)�OD~9�%�#EX#�R3,"ܮ�X#Ý��l����	��~��_�*F����r������_�qZ-ܣ����Gٖy�XT���?���ǖ�;q�����W��z��գ���a��N�c�"5���X��dWV ��q�Yh�ـ��Ϟ]�_@���x�u�2|�2|Cώ��]8��sl�j>�|�'�|���ה�F��;�Z+�/� �C"�J�E�52�������Z���x!\D���K�j����b�6/�5Lkkf�펱n�����R���?6|�g��朓���6�p�j/<.]#�N"Ô�����e�Z��t��TL�
Ӌ�8�}xx�N?��w�����Ğw���c�r�*�~y�+�n"������`;~<�?���>s�&M���"xgHo�d@�K���Ѯ���6�o_�lct2L�� 'h��?�aUC�i2���TR��g������g2�{�N#�.���5*���"��ǧ��dx���U�Ӏ�E�`lT�6��Pl$2쭑a���yk����s:�5
�	HD`z	B�&a��?��b1u�<����R<����DYi�S�c�P�55�c)���n�mS	�q�pr!v�xc��������X���J�a[[�y����\��Άl�z���^(�}��[�T�!�閖� �w"�˸���Gl�>�!�nnn_?_TUW�܃�w�jډ=iǏ{������)X�pvPtj���3��Db��ϰ}��S�3�c���(,�0e�b|����dB���!}_;�d8F��h �K=��zUKl^�L�B�^�K��T�!FdT�p@���S�c��[�����#x�ޅ���8��	��F����X�j�wt��M;`26��?�G,�l<��Q�K�ob������>w7����a"L���1��Qն�Sf�����Ay]����O�.P����Ʀf�eb ��_���z�cj��p�	D�ԙ8w�z_���g/Sȶ`h������|Z:��74
��,����c������,[�C ￅ�����A�?��<����cTT3������;��1m�FD�Ta��x
b%.�jG���X��n�X���O8f.X�m?��K7�k�5E�,BbU��x/���J��z���s_�*�_��vL���Q���	;�	�������k���8��49z�v��j6�X��,<_�,���MF��!��G>�(>i�_�C+�N�Q�b,]mSڌ|�b�
�q�H̫����q�q;�]��x8O��ÄPL����5_�c�5.�}���f8{yS���Hz��AXl&�������t�yF�-�p��0���l��&��1����q尠p��O�Y�?b*݈i{Y0
�_���4	�#0$�k1���B��|��4�f�0'Ry#�34-��|=�H!ݬs]:Զ���!�߀A��HC���k�a�c��?YޔA����"�QhU�sL͂���I0�z���%�т�*�bS�||씈�9�⿛3���ω�(>	����(֊���'�T���Ih���kn����o�0SB,2,�E���q`��y�g��J���x�&�n�u�=�����~=�:���'q��a�8����p��V�����v���VM$lcxnb�(�e�?��1�oA��GQ���W� .3q>�#�،T=ULJǹÛ���\=�7�m�U��ckp��8��*��zmY�������S�a�l�c��O���)�,����懜��;,��ci*���v�p;e����������8�w���r�%.�,r�^���Q�PI����8���2�[\��֭�ν{���p���ב����s�����0��&�3�^�x�έ�FZY!R'e`ˮ����e�<�����)×���5�����z~;vm_�M��`ǖ��t� �ѿ-ê�e�y�F�����`��w�E;e�ٓ�裌�^R5�C}�p���HIM�Xgwx'�+,���׆�¹�˝�>��ؤ�D�t���t�b�4�w����~�
X��#���8u�޹�g����K�{��r���]]Oq��mܹw��=�γ�g�WN.>20�����=>D�K�3��s�O���VXD7�,��]=��fx�kd�Y��>{E��)�W2�M?�Z���xJ�t2��Hs�?����[Q�uBl'bנ�A//ЉKW]ҧ��4��e�"�S|�s5��R�eX$�]f��B�c���G���%
:��}{?z���/�ڸ�S;X;���b���$�g�i��-(�v��������7J���+&Lp���3E��Kv?�.Npg�6މ����(��n�U��<�,-�l�jgJ4�Y�'-��RmGY�y4Rm�R77���Xʰ�%���'g�q015�{�������������9"08aHJI���/�����O	O�P��!*:</FF�m��ǧ�jwL�����F�x�pl8,'�cl`	�(���K�@���h��:UXk1��UT�z�N�Lh�8]�1�3F�[�T�0��F~�,�[�0yJ+����ſ�o�5Zg/�87/�X���ڋ/(�f�0w������|y`���ܻ�j��/�}�^xL��'F�`�CJ�G����l<��.냕���g=�x�:(�;�¸	����G����}����h�v<�㓱z�fU3IGT�.�b�}���y�!���?�'�����fӷJ�z_��;(�K)�00�DaIΜ>�q���|�t�?³�v�VT)6�h��7�~`l���*\�ێ��߱j�f蛏�6�@��QI��x�!e���ُ��x|j� ���cǣ��n�A7�����~�m��Զ��}mj���̧�_����`�u��k���3FY�#��
�Y�u2����!�|� ^��'�ަ`��7l�a�#ݥ%Ao��;fb�k��Lj�t�'�����W5g�<��{P�҂Q��0������M����<�Ĳ�`Faз���oEG�0���Ԓ�X���������Cs�\��������rj�;�#a<A�5M���?�?���L�E����v�tM7gޙ�n�&����[>��
i6�E<�4|��`R��FMu���jr����܇�ݾ��G1>|3�����ia��+5��Г�x���\�+(��@j˵5���H�%�j�G?��9��}��	�Sv���@'�odX^t�f��BA/��������Z�է
PH��=s�7�h|26�n�p�W{Ԗ�c��طk=����?��]X4�	�~p�� K������"�:X���J0:�B#��L��?zA5Dޱ��V���t���5e���
���ؿc5_ۇ���M�����)ëp��Z\:�Gv,��ĉ]�p��ho�'��?�;=E��v�q�z9�!%�!e�!�G�bbJ�U�
]Wk����[�����y�0N��mƙC_�ܡ�q��&�=��nZ���b�EEa\j6��+`�W	��j,��K�9t?�ߏ;���_~W]�S�)�"�Z	���LB����O3��w�p�W���b��V!��a)qX��3\�~���]O�a��~���=1��$~�BA�'�~�[�ۯ���Mxr�~~N�b���zN!ֈ𰤪��H'}�I�ݔ�n�vq�0��!�\C߽����~�w]�(_�|w�s�ט��{W/�ecbt.&&�#�`��nDb��J��0�2�$�� ��;R�u2,5������5�P�����(-�����hjkŔ֩(���g+�⧓�p��U|�c+�.^��m�2�5�����sGx�`Ǿ�z���=Dٔ�����?E�)������U��BH9���F��
�a�:�r,P@���D<牟�븖�8�S�U�XR���+%��5F�K�#���4p[<f+��U�F��9�t\��Ό�1�f��'2\
��z��T2�͠g�L^܊����(SRÔI�ef��\d��?V���m��|�78�Y"��R8o2L|�a��qa�a���eaB`4���UP���2x�G�Ή��x/x�!( ���@\L4�RS(�q�/ʅ 8�A�>� ����?/��x��g��\�ˌ�/��])��������{so��M�ĉ��@�O�O���t��M��V/�ys���GHX0"�#(������� F�0�4�hC=���(�_��)���� l���(C[|�o�1&00�`D%bbP2>Գ�������)_z�0���]$l(6�yp�n�_�l���P/sZ�~4�4��Z�7�3}C"_�2�����,�c|�KuM`�B�S�����uq�@xf9N�x���� -��ə���]���ST�5cźM��+���qAm��D8{������s'�_��s�>����z���N��ol=�a7����F[���; �Sg`��[�c�A��}GN )+�v�`1�	����,|�r-��g�}����|C�S`DE�
m[�R��:���������8y�2�}�^~A�x�\�=�n�t<y��?�ByQ֬\����C�0OSk�9z����.A��0ʨr�p������r�&X:�`��->ҷFPT:囅w�띻�˱��#}�y���E������,�q9c
�|C#Q����?��W���B}��U�Z������7%<���#��
[�����س�[�xяk7� 4:�}�@�y&�`BF��)ğx&MW^�H[Za�����l�)���lY�=���)�f΀��	0���OM�Q�:W﷫�r��=�����6\d802�fN��+b��7mٯz�����e[)>0��(�|`��l��Ѹ8���N1-��ҙ��S2����]��Q�� ]���{.	��J?�
N�_N��#��뻿���>����U����
rX�"�i�� ky�#���h�aN������[����=��Mu���x��N�^-��7i���=ʯ�D��7�Y�`�4��.
� �����u����$�����"��W��_)ǣ}�TaLP%�VĒr;B�?}#�"�Q�D~�L���Kt�# �s� �z��3�]���2�����xz��/���rPS_�iӧ���
�!p����3g?XML�[�d8%7��y�'�Ŕ�*�3?���o�b��B�����Jʾ4�(e���1�Q�t�=l�	n�ظj.�����õ_Q��2^�+G��܁��y�j��}-N���w����=tSn���tQ��=iG;�X#��c<�����`�'D>��"��,2|���E��;x5Ё'���'����o)���ԁ58sp%.s߮�߃�k"�(�q�p̘��հg�YՀ�[��ľÇp��#�z���A
-ً���2��Oe�����3��B�+e�)e���13��A���KdT� ����H���I5U�u���A�;���W���E�U�u0�v
������8.�߉��7�0/̙��G���o�࿿�kJ�+��� ^����cp��L��u�y�3n���?Ëv^�kg��ݫ��k���@�p��Ed�P�l������|$��'�1����3,�~	�]��)pL��(EDx��
� 2����+A�YM�v�&���v�'x�2:���EĒB��[+�QF�+�P8����г���-%�܂�9L�(XA�q�v́ر�X8���%��1!����lÂ�+��'��X
�]�4�Ƽ�M,�Qj�R;,"�'P�m(�o�`kA[ClE,UJ����ฮI�����4/�q}��D�[R�-�s_��Gb3�S�*��;c�8�����+���ɰ��2��&Y0Σ$O�uX����%��2Tj(�r��?CɰI@&�3a�N�4P�}a81&>	0�k�(�N����H�y�Ô��[��# ,����Edp(ғ�������xD��"<8�i"EL�8��H
ft"��?�bޒ�Fy��@w���">!!��c�?*!����/���p<��7���,�qQ���D~Qr󐝟� ?8�wd�oGX���=k|<��d�1f����xl �)+�0u��d|0�<�`�E��a��t����9���-���d�Gx�b��Eԫ&Ƒ�0���R�k�dUp��U�"r2�Vo��񛄏Y@~��~䖤�4��v"<�2q��}�~���$��a�����9z�þ�OQ�6�>|�n܆QV�$��'6c]������·�~��!&6��+�HXy�v��8.�46�ҿ��b�1�*�zЎ{O��q��E�v��.���w���w<�{����m��#%� v"]�an+_�sE]���'�<z���Wo�Ŷ�ߣ��N�.�'v�0c�,<�wO�Gs}<]��j�btv��z�5�-�Ԙ�mhޣ��_�(+���,�ţ���c���1��]�-��Kq��#<��w�;4�����B(�H�)��wT7�O�Q}�;�{����<�ǝ}�b0q������P��
Wo�?V�p�%kף��Ճ�'�/�d0��<+^v���pd6�_1Ƨ�a0�r���])9���=*H����2E:޳�h�@4��w��)���<�]�x�|`b7��;���Aנj|��)����҆��=e�4]����FY�}b4l}��'�X�qn?BV�4|j3���B�瞀O�KO�D��n�(u���=!��G�[��P~E���R�A󢛎�"�Vh�%�B��t��噾����(��T���-B�R���;���[Dne�%�2���q�%����0�z4�|+�o��J7n�S~�ʀ�/"�(�'�9M�v���v"��d�?l#U�Ct5�"+��2�1�j���Ū������g����K�	���j
&�vD�j�%�7�)����|yN�l'ݩ)��q�y8>F��2_�S���`�%M}���-�ϝ܃��G�p	&�Aa�d�����9�X�sa��W��^�>�z�?J� �a�˗���Ȱ>1f~)������O)�f�`!��X[��,'���W�֩͸~r5��\A!����͓����58�s-���������1t�.)�=�N�j����y�#Ռ�L~B�i��-nLi~�L;�le�ٓ{�y� ����y�}\>s?�یS��?}�3������8G>rb'&�j�gf�*��*�ZT��z�Y��{�w?���Oǳ�.:���H�0W������dx$�a
�F���n���VQ�K�RY���"$��+�����|����::ۯ�����s�eX8���3��0.����������+g0��N��I|B�~g6���4ч�ý<=�������)z����v��D�x��"���|�a��~�����X���n����8$������:ė-��{nbƦ��ʚ��F8P�ƥ�s3)�"�)��p@V3����{�GPR,������	V��o�k{k���A	��X;|dbkW���7��_��۱�jӎ��}���nGq�bxP�ܓ�*b�
�䙰O���	�)�b2vRkl?�-	�Śt��T��#��rJ\).#���t�l� �����G����geX�
'���&�0�c��	3<��Q�e�4��Q尉,S�����&�9�����,��^��aa
�1��)�#d��/�2��D�P�(��q��)�0y���-��p��A@4��hQ��b������tDFF�^��&�'"--�))HH�'q�O�AlB$b����X
2IJ�A\R"cBo޿ƫ�֤�70$>����<}���� ?xJ @�m�-02L����IY�MM�@&���|&a1��v^0�	�}#�;DR��a��0�q
�	3uc�(�PM�i�w,L�X 0c��)� [����'m.�y�X���,\�	O�ID���a� �P�bf����0W+!��8���<�A�O:����>��-<G)ç��U/}IO
Q��8K	����w���[������Ϡ'�C����	~��W_}���1��S���q�"�6s!�=Ca7!N~�pMG|n%������x���r���]?����ԅ�6s�,Z��w����%.p�6mم��|E�3Ȱ����f��}0����|�>�=�ƥ�����m(�����������Cqi.]���/^1����梱�'�UAgWV~���G��d�򺘹��=,�Z�"���?B/��;6����ܾ����p��3�Sh8�3���1�������y!�˞�v��K�j�Q2�3-��W��"|�I'v�=���)�����xM�[��51���Ρ�x�:�f4���W.ï�����G(,m��S L�CՇE�P�?r��4�h�	L̀|Mᛩ��5�79Dc�y J�
��, [?�Of� �	��s���U���z!Yj���)�c�~�vt��~ԣ�I�Gv���5~d����B����>�״�/F��#O��V�r$b%}4�K����P�^ ��kq��ᝆ��=>��ˋ�j�ZU�&5�)�Pjh���ÿK�Z���u�:�wgꖪIeo�r�b� ��C�0����?��-�a��[��߸U��s��e�v�:E��ȱ������ C༎\��4Y��������r8'��9�^�K /ך�u���1"�a��O��d>��V�����Ҋ�F��F��K�����a�k>��$9H��:(�~\��b|2!_u�� M��]Pe7	c�D����#�n��fpm31��&�KaQ���[@��B���H��[F�e�h�iBh�
�!�1	����S�s���ϋ�G,�a`e�2&{��G��S8�#E������u��3[pf�8�k.RR�؉�G����E?y�>�=�O�E:�c"/�=y�O�'�(�"��]Ip;�=~���jD�E��=��>{t7ExN�g�?o��cq��flܾ�UEpLN�SN�'�½����иb5~8|{����7 -Ջ��$Bdxp��o�ai*1R����Ι���r�77"��Q��W_�Ͽ���]x�� �na��]��<A�҆w��*�]���'q���q��:�=��=^�R���>����Pw��p����{��1�s�n��#iq�w�:� �Ƀ����F Ǒ�N����h�E��?��y��K�Ǆ�j�ԮDt�8��clL���Q��,8���Hq*e8e*l�D�[���;w��E�Fx�%1��I�	GBZ�S�D	���p�H���2��r	�9����������(ßQ����� �T�pRo�p��%R��H�EU�t�S&5�X�s����? �t�b��u������u:"�܎B+�&�:��2�k"a5B��R�-�I��1�Oǧ��O�5*`�]��R
p!EX'�٪��ѥrU*�,b,"l�V��E��'S�aL)�O6�25cj���a 5�~���L�����?^����D�%�/8n^~*mn���{���?��m��n�W�b×d#�ظ��z����}��ބ�L��X�EKc�9��`��Z��k�`�ʕX�t)._���aٺ�X��,]��V����KU����k��
[mo߿ŵ�1��.ΰ��[��p�����,ح)%֔��i�]�G)�'<?V<_V��ϡ�_1,�+aÌ�>���'	�"��<��a�0o�7�M� ���(�F�!6	��yd�B�؈�h�M�I�$�����7�S�p����r+Bx���"�:1�s�(��;:�����_��[`?Qjl8_D<)�-mm�������k�\�x�I�CGN"5����p�EE�2�8|[�EaU#B��G	v�
���,�|#�����Ǫ�Wj��vb�CȞT�	�'_{g��T6 ��Y�u9y�_ʋd�QYעD{��>�;3�	DLB*
K*�y�<��Bw�s��������z�3�a�b����+�q��u�ټ)�����
�"X�� �t2�����e _|���hO�c]����3W�`�A�y�vJ~�]TO"���8xLχ�}�,^��)��V��G0��sd|
�'�s���2a"R�'��46�p w�����kt���7o^�ˡ��Cww/~:~;�ÒM�xM�T��b kY��RX2ﳌf�a!R(㳗��S==<7::0s�g�+s������ޡ��p%u�<z�%�7���&��|�7x��t�i�2�U3 ?K�)/���1o�j������(o��1�d+��x���LLU�1��I�>YP�A�ʿR���=BdC�y�h�,%��|5�p5mr�m���� T/~9�6��#YV��j֗Cr���]��}�۞"F�����y��0�6�������!�E��M�%������|(��.��i�5�}ֵ]V]����cDh�5����7�8�气�v��Ei_l\��L������f:ǿ+��GI�����thz�ТDX#���c�ȧi�b4exѴۭ���xk{up�b0=�0L���W8<à���!����'޻��e0*�QP􃫠,5�u0��ʯ�&�0�j�	1�4�0�K�B���7��>�܏��{%��;
���`�8K�ĽKGq��f�VXj�����Hwf[p��Z�޳W}M��ލ�����et=���������",}�K���v�p;eXS�D	�3�������t�£{gp��^���k��v�?��l�ţ[q���Է'�mì�s���I�H�KA5\��>��Ӱ�op���S'q��=0,_%�ގz��0��������x�����n\��/V!����)���������JOmî�bD��̾�ݷ��y�'I#ý�Σ��"�w_��k�kqO���ˇq���~�0/�5���_����P;^<�+�r�1�)˃���.�v�ut�?���g��^=���;���]��}����~���l�� l�T��+���[�q1�a]���uL�t*�ȰS�,�l�)�Y}�,�2���]<��o��<�}����#�'U�/=u{�S��t�8������!�;r�w���}����8p�v��{���î~��剫QX��Y ���"��
���fX�Ԏ�}�,8������)�oh#����:8_�����G0V���XA���X�	g�9gJ�ݿ@I�̧�m���[�aD{a����dx�>��B$W����&����S��]�g1���+B�`�E�͂D�5M$4B���M�2�J3
ʱ�JM)�f�ܟH�6�/h����S�P���/�>�p�g�0��	�d����㼃�<g	�^��C��������o>�ĵ���OWy�
�<��X����7�������މ[�̯=|��̔�=�2�ʓ'���ңG8M�9wﾚv�Y'��w�������e�6���������K�&d�֧ ��Ű����χM�$��6d�BIX!�`�iĆX3 �
��eH�FNk�]L+,§y�s*�#�(�S`�i&�H����:ՆX�PG6��Gת�4Rj���(`�Ϡ%����Q��:���M��X���KGW8�\NA���T%X]�q+��G��+��Q�(*��c���|��j���t�"����q{7��k8�`q���]���
�t���L��w <}C���Ebպ�U3�+7*���£g�X�z#�B�U����88�x!*>���������w�C�b�گ���	�\���|;����c�a�l�n/��~:�c���������}._��\����u�!���;�OϨBX�#�����D��CX�f)����#0���{��_|�]/~�m��S`��g�^�	��6�o>���>����>J��Ǖ;P��J	�����C��4"&I��}?�#g�ݱ����Y�pGϝc�x�ǳ��������'���E�N�>�%i�oY�rX�V(�8��*06�6n)�/Ħ�������|���L81�r�F`L*6l��ōG���:V}[�	X�I^�{�{O��������I�����8�\������|���f���6�Qp�υ��܇��ӔC8����V�E7l0J�>1`^d���WH�����B�I��Fo��\���	àB��P�`�kҐB+&���i0
�"��7\���Ā딞+��,����`��/�	�5�a�T�^.�o�>�#�XH��&�Z�=�7�~�'_�咧{eS��1�y�Y`��|���ڌKO�ㅁ�,�c�f*��v��l�7�ۭ�y�T�iHVݓQ��ȋpLU�`�y�n�F �"�oeX�0p}7"���Y@)��/�28���{����=�RP}�])+���<�!��eN�
��Z%�"����]ʰN���I�x�y	S�N�el,���G60 l��Ѩ>\4������_�]`j�ܜ,�b�{��A�<�7Nn��S�n��3_Q������#_����stn�.��ǷΣ��5:�}�P��Q�;)�]��R�Iִ-~�.Jpǻ�ܧߢ��T.w���>�G��Ù��q��\<�7N��؍���?~���:LHτKn�ʛ�U��I(�9_��?�8��W��S�#1��[�_dX'��[e�W
����^Qn����2����ߢ���3g o�l�6�"��qe5(k���gϠ��0�������X>��⮧g��.�1�K��O(_�<��wO���������n2�0�y�Ϯc���:.c��9�?<��''0��4�?:�އW��@z=Ʒ_mEHt
�2b�M,�GB|���5�abe8�~٭�NoQM�'6�/��� ;�͆C�,��9J��0J�gO�W������_��K����m���/!�{�Rj�կ�0�^��x�R3,���x�t��r\}�����Ȫ��	Qep��p�)��Iӕ��%j�O�M	�C	f�Ly���0����B�ա�a{��������X.?VK��LU{�AS+m�_@I��f[��k�+�u�4J�T�&��pr3�bI�`�3df��ڮ���)�Q�,"�a&]1�6aa#m���Rf���-�(�a��,$��`ʢ@�q��\���f!9���0���\���@��a�3�lX��:8V����fs��M��k <�ґW7-�֢u�L�l�.\�)s>G��eh��9�-ZCV����
���3�}�;�a��/�8g1���A������ u��v���^���s���B	����s1y�B��٬�=S���6�i�
�5� ���	0pu����5vep���;;i�T��,a^��A�ꪉ���E��\����J�o��f�1�YH4Q~[x��3o�i�|t��ҫ�a��R���p�p�d�Q��c�Tj���,��BT�O<�XЅ㽱>H(k��0�&�$����&��`l���l9{U������P�M�O$^��*��/��c�ӝ��QWW	#���LOť�W���.�Ee�"&N���������s��Qb+݈y����d2;��ת����׸�����o?�
����|�Ś��W�Ͻ���W�S؇Wb�}�~�̘���r��`��ոx���iGc�|x��7$^�������l�\�ڻ��3����]H�*�X�(����!�im�tn���kJ�W~�6҇��'�C1��ye͸�����]�H΄��7��y�!��@�-�MB�G<�y� ���	KV�EiU=��S���u�8~�N]���+�7a���)�B(כ[V�j{~�����?���"$>^�����Iȇq>�Ja���j+Um*㟭УX�N̄�C4'��؀���8{���/������,T���G7N�g��2��t�~�w�w�{O��QP�O�l`j3��0��ǢU�0��/���e--x��
������Q��a���}��=���t����Q#��������k{fx�Cç��Zb���t���9��'>o��B$����%���>�E"�m��>ϟ^ �%�1���Q��@1ףh�1Fs=����l�S?!�Ӹ}��f*��ש�nc�?���7�Ӝ��+}��@��ꩾ�u�S
�/n�+�y�TvC��K����Q��c\��I�g~��ڔ����1��1�u<�ZK-�U#ƪ�X$Yd7�]�}�F��4�S��6y�Mjp��gi�˄F��H��R�[�Fe�GJEǭ��Y�T10����b��0z*�BԸ������X�5��c9�6�3�b<�C�g��<R��]|X&GT�@��O�A)���ya�����.����;p��7��/US���V����q��Z�>�	���2��2|����g���z����	�ڟ��ς���
iR�����Mt<�����q��^�;�N݀�'6���p����6�9�w���=���ꥈ).�{�$��@h�\׵!��3�X���+�~�ާ�Z��?��?+�/^�P��j�������5��5�~{��]�{�$�~���� ��93>C�Y�Č����e���%J�P'z(�=Z�a\��y<{L�}|�'\�O\�_�`�U�H/ޮk���?�2O/R~/
�����||�1=��vJq���>�wc��m��~�F��#:��H�@p��W.���f��M�Ov�3Z�6n)��a�O�b�6�"<[�9Oӻȇ7�OZ?ێ]Go��������'8z�Np��S�p��U-Wpp�N^���p��e9s'.���K���Y��<�9����A\#��*x�t	"�"�Q
����[%�:	F�k�����i
{J�=%S�n������ZQ��
:ɟI�?C�'����`�����Zaۤ&�è9N2�5,�!EM�z���M�	e�,�f�R+Q�̧�b�O��B	,�)�D�K-qx>,#
`9	�QE��.V�U$�:L�`�zHH3�|�	eXj��� �ܦEh6�(��O�#�w\TƆ���7�.�0q��o"l��`�3�H��Dʳk8,��H(	�@X��5$	a��pK�x��'�����}4��2��>0t񂁋'􈁛�b�x�yPr�T�Q�C��8�v��A�@�w����p�o�S|3�ê)�e<�r7�V�W�,�DU�4�&�0����I�4-��MG�Vҩ,�Rl�y�(ņ"Ŕh��;��AdL��a��e�9\K&���db�}bv5V��K�����1T7πG@8\}ào��is�G�����vWR�������މ���^Y���H��Ł�T0�������Y+7c�ڝ8}�Ѩ~�`��r�l،���R"���W��Fjm>��]�JP<�U���k GN���kwUM�+鎍� �h���o?x��?h��1��O���ڹ�=G�!"1��a��	C7X8���Kl�s]�*�޺� rK�`��Om`��Q����"|��[��z�_�w�ry�ep����;F���3�w�Ń��������1�&|�� �>F/�㞣g�d�&>���<��ǳ��z�sWnb����On�z�N���?�{d&�j녿X{�c{o�;L@V�d�g�m�{1o�8xE�?���C��Lz��6��0����o�t�e��g%�^1(�o�O�.�No�?�)���y�m����P�_c˞C�Hʄ��bSr��O�0��z�=���.>���x",6{�R�c�|��W��CP ��	��ɕ���bH����{$�G$%�x�OxO��%Q�G�O֒�%UK��������u�\/�ʿy%�}/nO��o����up�t��x�3�������jIyӣ��W��f�W�+�Tu,܎�@!��4m�ߗ�&\���&m�Ӵ}��ZO`p�E�W�����q^=
��c�ܵ��'�p���5*ĸ�zT#�Ҵ�P>�A!����H1-�"�kj�G�R��|�CD��/�zq.x2���ZHא�R#i�@15��S�G��0���(��G1�ԓf�?-ëX�Ԩ6��`��60_-2�j�e_k�?J�kS ='�K���s�3�8l7�"\K捶�SX.�0ߤ\s��!�`���d�1�źU�p��<���Oo�
��9|��J\;�׏�#k�F�:�-Eu7�_:�G7O�ك��{z����ߡ�Š�τ��{r��_Ó;����qܡx_<������r�B|��7�pt+�ݏK�wc��1��	!���a��W;��s�0y3g�˽����8u�,>~�$W'�#��������^��o����������� ��`���N!Nk���K��4Q�H�iE\I-��k�S�ՋsBϳ3����q���q��F��F��xF�w�ǫޫ<�燧�G�?<��Gg0��,^>>��N������8��:t��֋��AAE�D�-<��R��I�J�K�Qz��7&fM�gz<��(��9}&�wo�y�ǹpH����p�$�qF�������@Z�dV�Cr�t���BbQ+2*� ���ӐP8�� qRI=�
ꐘ7�i�
k�]ֈ��F��">� �iو�*Cx�;��[�8�(�I3)��t
�}���8��t�FZ�|��]����|"�:D�55��V��x���+~��A	��[󁷦ۈ3(����53;�DF�񔧨J�W)L#J([�0�4��F�q��Bf�^A�W8|3&�A&��lU��b�Ɩ`l|9*�V�.���Ka+�F�_�1e����%�-��}k%�4cX�R��"�a�	[J�Mx�C3`�k�4�p�&,X Y���e����i,��=a�O���5�.��[�8S��\�{8��C(��	���
+J��,$����`��x���6,f~�s�� y���+�!1��h�Č�ᩰb�l&=<��܆izzP0C7��ۤ�#��H(�F̜�(�F�a�L>�����������6��P��(�L�e<B2�fN�H#�Y��FK-���D���~o�-�B=��,Z��P=�<��<�Ɨ;T�7�#�2<�N�X��v����3H�ƒ-���������=8���.l��&z�#,$?�ً!�.�`���T�X���kp���~JA�D��WJ��Xdvۮ}H�)����C���kQTQ��wq��/���|�eR,兹g�/�X�V7b�񴇙4瑚�J�ͧ�1g�Fظ������a�vFjq#~<q����y�Kv�=Ǟ��"���	�!;���1f<�|�W�����/x�����G/�C^9e��Ξ�c6ɹ��{�8z^�F�����?#�����(�iAVY�����7�aΊ�������X>���^a��ox����x�,)�2����MbY��t���X~��[�q�n'f��.�s7�pL���-���$�Q�Y���׵�l�:�5(R}���;���W���_{܍:�i�{��U/FQ��,Y���/�Iϰr�,��k��~�.��]�9�>�w{R�;���y~��W��P�xL|���7F#���'$P�(����[�Fޟ8�DN������~�c������m��ѥ�
<~�v��� A�Ii���[DTy�)��Q�� ����}�}���0y�#��eB��
�V�e��Mn�o����|4�rK���o�GdYɹ���v҆�
����W#�\^����\R�W&>� ��%	�Ty6>�~���R��9�W�L��a�V�b��F��g�)�"�#�+���Q��Pv�8�'�d5.�w�
u$���I��1�2����f|�m}�y>��Oc���z�Q�ENfySs.+r�ʼ.v���QaS���� ʲqD�4
ql��&%���.A�Im�%�iEl9.�FHs�H	��\��g��'n^>H����M+q��.��N\�i���2��|�kG�R�W�ֱ��q�K�����<���.�����t��w�{��ܿ��6:�^��[g���1<�~WNl��#�q�䗸|v.�ل'6����:��wo���Ӑ����������l���isѴf%�\=���O�������VM#��F�_Q���W�B����dF���s�q�VmD��eȜ2��g�p�
D�4!���׬ǡ��p��It�B��M<�<�g]�y���r�^v��K��K������{p��O�ey�)���Q�3���'���^?;�_������MA���6vڍIu5��M�sD"\c�RЂ �pt�"Q�}
gc|z<sg�#s&&�π{�L����¸TMͰc�8�2�5.�0!k�z��!�N������q��+�mH)o�b8FV��v�
my�چP��I>�7JIP�)I���ĸ���ʅ{\>�C�168����L��FQ����qSG�Ҕ�J��S)ǔ�wdX�s�R������`��A� Ɍ@����b
��!ќB'�Z!��P�u؉Sx�e��F�m����BX�'3CHl$S`��;�[�����@SN�#���P�#�8��0��3
��@�5����Kʰ絎)�M,�7�LI��aU�T�I,EXQ����ܦ�Xd\�wD.LC�`�B=@�2^`:̂��{��~Y��Z K��9�?
`/�pC�y��q��HH�\�G�$6!�0􊃞G�'��*8&~�0��Sݚ���?�!I$Va�pN�Ǆ���T�a}�H5��O�&�CB$��� -�x\D�D��D�0eW�񪶼Z"4E2����*)���̘)��A8���HS�(���k�a�a��+!n�,7Q��`FL�)�1��6t5<��o�躥����n9���Nc��c�gfc�sL=�h�ᯖ�p�*@Ɍ5|�����?Jf���}g�b�O��~�ۆ��ٰud��)�>Ǧ�c���X����m�g|1,�c_2s�n��#���|��1�ܲ3W}���������*L[�-�"��1��PB߀��~Ɩ���y�,�j��>C��/�h�n����#K�c����r�~8{��Gۚ��ea�3�8��L'&!���﹀=��a��{8x�G�ub�g�|��;&�����Aˊm�q��]��#7���;�BiN�񘸆�9X����'%��+���]����>�;� k���m�-�sp"Z�o�ԥ�����5e�>�8�='o᧋�����]�n�wG����o��aH��lX��g����W���=��q^�x�ϷbN	�q��DpA	0�=m���40���D���E^^����� w��%s�V`�˸�מ��̭'���Qd���qEDr>v�?�{�x���P=��MI���W������?S�����n�����0n����0�9~nI�q>��d|D��H�8��c������?�K�'#��A�G�@:���/����1@��/K�	�O�r8��lM*��G�Y�X����
y����a�|�@�ߑd���!�{nO�Cr��h���%�d*>��7L���R�C���;%{$�=9?��|�!pߵ|�q��4�?���7�vm��xKO����g�͂'a\B\3�+GM�[#WJ�eX}RY+�cB�/S�PJ��؊Z~#�d}J�>ףDX�F���i0�k�^d=>���EP����jK�e�jAٕ&�\�q��k���)�2�<7���{5,S�v���L���3��d>k[�2�"L����0��5��7e�\ G�=�a)p���D_4�NƖ��p��n�8�.Sx/^�����֩�����8�׎o��7��o����h�~ �׎�ɕS�4�\=��~p��_:����K?�֥CL������͸~�+�9��|�����S�q���;�?ۍ�떠��aYY�-�Bl�|�Զ!������;?���3����>��H�`*�����_�a�4���W���5^��Z�K'Ȍ�>{�>ߊI͋�Z;ymˑ޲q��S7eKfa�O�q��E<yyO�/�����<������Q�J����q��~�����S�{�I��}�uǯ=���~���?�ǰ���o��DFM9��#�� ߼
�LAX��L�U��]0��[��{�l�ǵ[&�7c.y.�(�Na��yd.���K�<����s0!���́{.�Y�i�0!g1Y��ًnY��.?��z���Yp�j���iL��#��p�k�[^i�k6˘�[�L�ϰSJ+E]^�	��*�6�#i�|(d\�9m�?�1�E�@��GF
�N��B�����������(k��Bm��(�o�U"<B��?o�[;��X�I�l�)K1���2RB+�L�,��JLc8.PvM��B�`s��S�[r9�4�[�piz�O
`"Ôm�J���4�'Q�0�N��0�mrA��I�Ƿ��޶��iҞ�0 F\�q�S�5�7N�L�`(r���Lf��L�a����l�P���xo�)�K(��U�x�E*|�'}3 sK�AX�|��O��d��K��j*��y	3x#N��af�J���a3vJ�a�4f�a
�`�iښ�w�X�k�M3�j�u�y��y�`N,X�X� �bjKI��m��b,ESJ����5,8y�Ð1@����R��j��^q�Z|^/S�{S�L����z�$TbB�d�1��k/A��{=���2(�B@^=<�*a�J��dxf�܏�TP9�*4j��;O��3��� 0�r� ��גA�y@�y,y-���݀@ʮs�d���qKZ�}vd�娐2�m�\������Z�����͚
3ʍU`ly��Q������Q���鈭Z��>Y��i0���y����"K&�0Ȓ4�d*j�#(���-�T�Mv�<������7�)�i��P��9H�Y��I�aVʠ-K��o�k�g�7��^%R�עt�Nė.A�̍����ES�����&(��(�����m`��&@����c`l|�1��6��*��.D�/P>u>���a��SGx����z:�,�s�~�y+�`�g_c�]��t3�2'#<�Ͳo0}�V��ނ�5[0m�����K��c#��s���F���1累E`�)���>e�i�[>�u�$���>� �y�$����׶�e��	������������	�F�L���2�1����y?�/x��o�$0��c0I1�0��n�E�v?	��?�n_G��",m�?���D�����sY��tD)�b'�.Nz]��f��F�� �3�Ʉj6!���I�1�a��j���<B��%�`)�=�M�_s�_�U��u�׊�YG7h�X!�j�U4�2
�4yP��gjS�����2<�8�#�V�k�1����X��u:�6�9�e|B+�Ʊ,���F0�b��[��2�2����:|�un^8�'Q����#;q��f\9�WO��p��8�w�>>�	������?�����w~/�ۃ[gv����pEj��^<�.s���yb+��O~&G6���s~7�_܇#'wc��U�j�B`eB��8�Ms�Pߌ�iS�p�r�xv��:���b�y��1�ׯ���Vz��?�W��k
�+�b"�Ҏx����|���_B��(i[���e�h^ʃ\���3]S��EӰx��yb.�?ɨ�2^���^�`�==��'g��<��^w]ī�x�s����
���e�"^^����hﺊ��b٦ϑ[_ߴ�(�pK˃ߤZ����)�՟��h��E�g*!�ț�ܹ�ș�p���fIM0�؅��Ji�u˦@"ѹ"�\&g>�z!�+>S��,"��H���fʋy3(�31!o�X��șAڸ�����K�B�OC��J��*��qj�HZ5�O#S��qi-op$�*ĺ�ci^�����Pd��k��92��6ȭ�PxGb�x$#d��r���v�Md
�|�dfJ0�)cZ
Ӹ2�ŗj�+�9S�-�Xj��-e�S�����!2n��,bJF�uH�p4�O�6��dS�L����B�P�LB(�ҶX�K7���8X󒟡��?�a�.����8�f�{�QH6%8F��_!��a�H���"v�2V�E���x60�-P����a�N�JS�������y�$��:��2\��z2����iLֽ(�eX��iM�YK��8����䏨�`�EI�i��X�7�A�y,a��)��J^$,|�Cʹ.J<	� �Sz�Y��^6�Qu<�)���zec^��r
(���eG�lªa\��X��!���M-��I%�y�K�ٰ
�g�S��r8JO4,���_㸯�,v`�g�m������2��}T�۲��]T�#cc�x�ym��O�tř��K�R�^b�ш�Q��B�?a���-�J�3F`��*LHg��{G������H�Chl�F� -幑�@D\�;�-�.��ў�|9İpM��z���<?�<oŰ/���n�kʈy�|ܦ6�<.b���N>���h�s�c�� ���O��x�}R06$c��`���QI�
o C#0.4
N�1p
!A�Z��g�*d\ד��D��r=i\_:�t�#��R�9-(�l��9��g�Qz��й�9/�c��7��ֿ�IKb�`@ ��I_�8)�c�c����TQ�Q�F���c�|<FQ�1�%�m�cF0����1�XP�bL0�.�(nC��a�v�孑p��R.�m�,��D�<�]�uHW��ѡ\����������HCȿ�>�Ub(�Gb�s���b4ɑ�I�RYQ�F+�SVQ�*3�d0/Az��3oҋ���XO�5��"���V�ày�A5��rƒ�q=F̓��	�o����a3�9#eX#�D�%/�<�J�����d��Z`�q^J�M|l`��Im�a�t,q ��?�t3�aN	^�_����+�k��"xR��Bb�������|�(�\>�G�Ǳ}p��F\<�������%��'6��M�}�[
.%��NN���NQ�ɥӻp��n��.5~���:��~ގ�����}�'��P�߶�_W���%H�ւ����<ym3���Jl?���5������;`ϕ�DxX	���XǠ��ߑ���KdX��V�e�寿�o���йk����.AV�b$�/De8����%H��@��f,ܸ{��ĝ�g�?p/����=�~~/zo�^#��㹼D�/�8�0yqä����?�s��a����S�ZV ��� ��~�5�Ԁ���<��W4fQ�g�w�l2�����d���x�ϧ(St)��y���+�:]+�3��j)�C�K��GD�5hDY#�dX�X���:�St3��V�ݲR�)�Y�5M3���Y�9��Li���jveX��S2[	�I��[���j$J�G�$�vE�Eƅ6U��d(9~[[���X�ɲ���%�i��5�"�-
�6�N�.�TN�gp���(�i��t��&��J"E.��"\��B"���9�H� �@�"�I�h�P
�d���a�>e���5nG��M��R�.�@q�-M�Oeo�I�+f�R�gQs��B����E��S�|~��e$3��"նٌf�B��bJ�1�r)�y0���>s��1.��ka��B�?�(¦�9�����zr�Q��>��4=oP�D�,(/�,Ḷj�^��N^����eX��Yh�afoK��ؚ�+���	i!��Z`U��.��N��P|��8���)��.���Hj�k8�����c� ��O�[qy���/2��v�qm��|5�4�OX%t&�fSjgQ��`�L��Xڲ ��ڱ���6��q�"��uL�BƧ6�1Q��da�c�e�"d~N�o��d>�ɳ�$�������6���烩C��x��S�=n?��"҉zU��g�ψ��v��g(���O�j�)�����`�P�e�mz^O�w6єR�-�[Q��"�0��c%������B�s�3�:��W��y�3�3���uNm��/+���aA��z��:��z��d�7n��ɼ�'�6�� �q�M<����j�3�i
��� �p��feYpMD���h�|-���Eâ�иh�����<o	Y��y����4�܄���  @߿�ߒl�c��������a�*���b������>�u��+��5	�a�X�c��{�8h2�E�$8�'��\�0
��1�/�
�;���S�<�7��B�����&��Q�F�h��E����0 ��2>�Tk��\ h> m��E����jJ�Qͼ:tp�./)�_���w���ȀϹ������M���Dr�ѿ���� �+����H��KyJS�G ӌ�Y��������^-�k&2L�5d>��|F����:��H��Z��VxM���B�Sڼ�ϥ	�2�e&��Ϙǘ��A;�$%��L�]p���7"�g��D�.�,$7�L�¼��q2%�ϿzބDJ0q���$2oJ���|�]��(ą�(BHZ.��0�u���gN���%���p����pz.���B�n��w�o���[)��p��v%��Eޅ�\���ݔ�(��s��q��n\?�7���5��n���ˇ�ծ��ׂ��j�oR[[�1c���F��y���Kl;rgn�����xH��B����b��9ӷ"���S~u�Q�� ��	����+	֊�n�5e�S:B~�]C�q���,Y���%Hk��ȊiH�6ѵM������J��T�f�T,Z���l��gq��e<|t���x":��ߎ��O��E'e�;o�꽳8q�v��V�B݌�N.DRq"�s���в��l�Y&�LCP�\ρo�,�N��ޓ(Ă���o�̛M�ɝ	���p�i�K�4�E�g5�f���Z�;q�i{G��l���N��1�HW), 3fQ�gRHex�QvU��9�F�)�y\w�����i�8�m#��o,�)�#�I�SF�I��2�Zg�}���&�>Y^�S픵ê ��d���-:�����R(�d,���k�x,�.}
�S�`�XM��Y"I*�9��"��ɕ��bM�Ia!)L�O��cZ��t�Zd܁�٧�K\���5�W�L�6�B�u�1#&�dl\���mś!Rb�a��BQ�F���q�p-j�H�집�B�#m���,���3�l�Aj��(�i�<�
E��c�D���BH�	�gK��Z�@��h3b�˕�`_K�To�,�<��[IU�3f��PPZ�~$NbMY��4pyS��)EU�/ȲĔ�����L���l��[py�	�����W��=Aw�H�{6��1�bA���h�����x��<��0��D�>J�Q�1����xn)Ea�
s[)�X`I{i���2V�g��J�`K	������J��+5R�
��o&S�)���C�No���Y�N�:������W��˧�m�r�E�)�)� ��e�d^�*����i�A^ �}dF901��"l(���Z�v��,<ǲ`�����Ky�������o��9Fk�&�\%Z���6-x���_9�\/�����>r�)�R�K�"��߾2�N^��1��7�<�ʠ�%�jπ�.j�b�x�!\�}�#���lGε��|G/.���J� ƕ����;�t��;��#�F�Y��}[�[��U,�U�[�\�k��J�12��D���:Vq3Ҏ�*~�U����a�{ǌA�>��P
UX+���)�[)��<��i"�L����؀"��M�S�L*�0�$�F��F5M�w��S�j��ZM#���ǴM��L�,�πK���&ՌKo��֐��P�PP���s�w>�6	�	���>���B�I$�c��7Tpz�>��`Lq6��l�+x}���9�{�6�yeX^��f��(�e� ��^�����2��`�q�_M ��uj�2�qS�w�f	�`J��ϫ�f�#2��B�*�i:�_*�i�����3Iɵg@���|F%�ub9�,X,��]'��GX�OgP���������N��v|�3����Yӱr�����8�0�^ډ�v����z��{vn�ށۧ��|��(��N�����uf/n�݇����
�K�xj/��\�aܼr�n��O��bͶ5��یԚR�Ϙ�ܙ3P�`�>[�̖6L[�v�|��Ɲ'�����=~�׃ai/��a��y+�CxA����6��DX�.�����A`��Ktʧ=�����_"�y>��� k�J��.A�����mEbu#R*k�^^�Iu�h]� �V���u�i�w�}�0v:������͏�����h[� �sZQ�4)e��.�@lQbK�]V���:�U� x���A����,��I�)�L��(�m�ȝ�� Px�
��.eW�י��,��YO9�#5�V3�iΙ����s��˛r�,Ι\GF3ő73o^��UbI��eonADYj�7�	fs�ӳ�j֙�mȾd4R��i��4���D���mj����a��v|xG��fߎ��`���:��NrDx�k�ZMz��bE!�N�� 7���%��M���ɰ�Y����;^?�as�%&Vf+F��h[.+��ޱ�,�����`2�CM� �>`CD�u"l#	�l�ܚSl��7Ք�HG�n\�mRa��dX����2,"<R�M)�R3,�+M$��R��-qT����jb�@�N(�h��r�B�Re�sG�����K)�"]����05����	e�$�Ô%�A2��%X 	�c��I<�rb6SnCxw��R�$ՠ�G�lj�G#`r�W� �׏�e��D�Yj��I����O��&^�V^�鰤��Qr(6&1SYj0���Sx,�f���q~��1�z���6�͸]��&�gSx\�q���h�}�Wp_L)�U3���<���}�+J�lǌ��f~M�	$���]pܒ�X�QI1�5�!��e���$�����(r��ו����'��f�mJ�6�y�!5~:�y+7F�!#�gI���x�r�c�h�Ԕ�M0�yV���wE#�^�3	�L�>cY����	E�T����ȿ#�q%(^�+������X��$�8p
���������El8x�Ӯ`��琿�k>�U�vP����'�\��t9Q�����_�RsKIգ�*����4���?��1�5s�V�f��t�N�Mal�谩�eG���m�1"���(9�uO%�N�EB%������6�zo�}��NjEb�D���0�39�����dV	��GS��V�5��u~�|��%�r�����@ɰ\sA'ÂFx��M3��+�\�-|n��#2}�|A��R�^=�q��-�H�L�+��K ��]$8��5�y[	���;�WS�&Z#>�B�4	6�tc"y�	RS�J����8l�@�2�ϭzv�G�a�9�K�V|�	�% ���O����<���o�T:��4�M���*��V�e��Qڔ�L��p�%���SH#���6�-���3�?�ny�?���S߂2O*V_.�R�����8|z�\ޅ�����{p�2e���}�{�9���]��9i/����sq��{��\;u WN��+'���ܽsWn���?c����a	Jf5 ��Y�M(Y�sP�Wb���[�܋��n�qw'ڟ�����܃�}�x����9�E��2,"��"�B+�"�/�(��	�g"���K��3�ա>��O����_���bx ����Wt���g1��M���r�oBڜHj��,F��%�m�$׶ ���5ȡ �NEq�t���Bi�L�N���i�1�y*2jky!K�UH�������LF����6"����_]�"�5/e��ų�U8>�fb"�ػ�B\Ъ�7��u�L�{�T�D��r������z��ԑZ-2\���﮹S8/Q/��r-
לf�Kv��fY�k�0U�4.��Ȱ,3>K�[�����H� ����j,�R�R�&�_*��U�3�/��2��WN�;�Z��Y�e�]+"����u��O6g�/ؖRa+r,/�i�I�Fr��R�b`����6-)I����\2���͑��1o
��7)��Q�'c)��)�X!�
�,L��oa��j�X��j�ך�!�NS�J&�q
�H� ��q�ci:��D��W��%���i6����i*!��-�r%b�Y��(�Nbᯑac��g��˦x�Q�(�հJ)�)�M��X��E0�:�	���ua�CI�����S�7����H�F2(M,�4"�V~MX8�Jmc�%��@D̈́�H��ی���7��ÂL7�y2b8o��Wq�D�Rkd,Dp=,��娀b%?R)���wlY������#�/�*�U�cӓ�����O)���Q,`?%�Dp��ba���1�l��ՈA�<C޷:��X�&S����|&��1����`��� a2�yn���H	��J�Oe,�+�ؚ�>S�|���7�2��@��J���f�@ƀ�+x��a}Ϋ�}�g����ŀR:��	eKMQ݈��1ZF��}9��`��hJ�,#]G��4A?�BG(	�C�#FL)��bʶ`�`��ϱ!eܐ"o �]��N_��E������">�E�Q�|T�RƠ�fB9�'>_
>S|��S������aV��s
���a|x��rM��P����0�˪���M�SL��H@�cR_#��"y�y�f��f��sB�My�߄1D�A��9�A�Փd-R��i��v���^�1\��\a2�V�g+��%�aA�>#5��������|�>dX���i��%B�� ���(��^s=>7��4�"�E��(��)�������B�N�!���rlB)��4B���2<a	ܭx���ٰ��si�"��0`3��j��՘��`"p\I��kn�q%��M�~*_C�����@%i�Jf0�Γ���ئ��.�M!/�;���i\����+p����o�����5[���N	�N�ս�Ĵ`&��2����Y8E͘P<%-�(�ǔ�a�����^� �E-�ր��&��4 ���U�ȞR���X��l��9�'O���?���}�C�^؇��S~5ܧ?��>�p���p��!\9uw��ã�7q���?~��mD��Q8���&�`~*W.A��e(\�K�a֦������~�(���}���4�~�7���%%��0B�_hj�u"����'��_�3��OeX����~�S���D��_^Q�#���t��`���9�
G/���M�Q�x+�nA��H��
��ܖE(�� M��YݢȨjAze3�*��Z1�H��GBE��T�"��)_E�'�MHnjC|�l�N]��i�M���� �v1�j>C�䅈�� ���V5����T�Fp�,��@@i�yS��N�o0��&��L!��Tƛ�W�L�{�T2�e�+��ď��-i�O�42�]��͘X��'L�D��>�Mj��&>M|�f>���yH�у�A����{�1z�OPQ�wʺ;E^���}�n~v�b0�RA~��k�9UE�o���һ��wSif2���y����h�a�lF�ܶ�q9<&q�������/�,���PȠc�|��ί�ٟ�L�-���t��Oo`�U��K�cF�@%���5G��8��,�ǧ2��4��;q'.�[΁��� G��8��K�&U����H�+I�m"eY���<&_	�Mb1l���A��!��gqYʅS~r&Þ�ͩ�53O��yJ%�*Xp�,T��q����aE���HA�0H�@��cE���Z1��b fŀ̊�m�s`�}6O��ȕ����gN45�Z(9���[��I^~�aN��Hm��ΒX����O�O�93�&��&�U�UjVP	�D �(�f<��O�y
W�;��2�(�3��ZF�a��iɄ�TΔ��sb��ʐ�c��2H"��~�c�`�m�i�;��Jϧσ�i�ke����6��s�����K��1�y����\�'P�&Q0�a�XJ�i���(��.��B�;�+�4k:%�A�>�:=
�Z�ǯO�����uӧ��ǷP�)w����T����P�b)v��z��zq2/ŗ�Qj��˨�ZDz)���6�n�5M�[��m����51�5���g ��k7��q4�є=��~��Ɩ�àt�- �����IQ�O)����"|8I�Qp!>��^�2b�b� Ƅ�5�y�`�#]-�0�3�=����1�Bh�B)Ua��0^� �<r��	�9�q�(��\��QQ�*������/i"�C�"�[A���/�u�H��1�Oj�Ǩ��A�A0P�*H�[^o-��=��� �:�w�:����#����]^-[��p��xL�r�R6y�o�-�H)�"�:)��m"��2��b�_+�&Z!���ل<�_��HL�2,�Y�'��6`�@n��J;_�p<�=j"��7��3��>��$
.�� ۥ̠�Π�Π�R��%�׊kC�M�<��aO2f�1s&�#i
I��+�d�iN)(֡�]R�s�ʰ��%"\(�\�GL���K�K��C|�ǘ���X�&֭�O�"��φ_m+j��،��$7�!���3�Ѷ�+6�������O�p���B��u��_<<��xp�^:������q�4N;���a�7_b���0y��5 �4�6%+���嘼z�W�E��n�Q\�������)�����!����}�x�q�`�	D�_R��N�_S|�!�俍���#&���y�A�_�"/)�/���^S�_b`�9��ÿ����øx�1�ۂ9k��o0c�zԴ�Cm�Ե�BC�lԷ�DM�tT6NEeaZVׄ��:��7��i*�j�SY��ɵ(��G!�$i�MiFa�T��"��M���i���4��L��܆�ȩoCV�4d�P�'7#�j
���TR���B�.�p�LFRq5���PX��I创T�X���E�+SR���*ĖU#��a�'��H�%�˿��ӄ�R��#4���E�)D0�T��M�	�/Q�� DK0	�-&�
�o̑OF�  ��B	�]��Vs�/�oz1|Ҋ���/�~�����o�U���P�y�J�_��|��O:י�[G��70�A�5��õ��:����I�H*0�����/�~y6Ȅ�ɤ�Ծ�}EF��3�V�3'�-��\�{F5<�&�3��9u�����r��S4L����=nw"���y��^�8i��+�>ٵ�/ޠ�fMjF � ��uz�s;�_ϴjRE*I��K�eB*�-�P��(]��Wʎ���K{Lr|2&�=�ZKǙf0�>	��<�
R��rk5���8���U�"�N��^�mBf%����ם2<!�� n<�ܶKj5%�$kp��	%�%����=���T�u�+�3븞Z�e	\'Ͽ��;SW��8J�%�)�Δva<��'�r��p�������U��0+(�Nę��Hyv�<�P ](���_WJ�%֙���1!���ܿ'<OPۄX��R��)Г(Ӆ,L1���� �1��p��A�=�<?�c�d8���tq�=��{���#�����\�}*�4����8��q�&���x<D���t�d�R��.�(c��al|)��q=����3��8���x�'�y��R��	����x�Μ����R��5� o��=��9tm��i�}i�~e2UH3������xlZ(����3��~���0���`�{�����kb�g���j�se��k������)S^��25n��Œ���c
)2%0g`!� �%�PjJ|�ST*a��`�uZ�7K�C��Ŕ�w�P�h)��	����T1�򏆪��RM�$�2gPdB�C)C)C)�#"�#�(sz��'��Q8�kdo����pJ�>�xA3n�a���b�E\Џ�r��e~�eД�)53d� �9�A4e:FR�������\��8�׀b��d
�6b`a����)�=�ʪ�.���X��F'�[A���K>̣�`�_�����sY���ZK�[�_#���4N��I��-��}h��`����fX�>�H���F����m�n�|�9�uF3lx��fOUȰu�L�`C�=��H��pΞ��wz��t��Fܳ5M1'���"��T�4��<y������zO����v�,�φo	)���y������X3�9M1��Kܰ��BH�*�5-Gx�b�7.@d�\�7�A�Y���HihAV��4�lz�ǜ�Wb�W_�˝۰�ؿ����O?�űc�q��O8z�v�ށ��6`�ꕘ��34̝�R=6*Φ�.B��%��fZW�����]��+�t�.�芽Ң`�",�(�tFᥖ2M���x5D�%R�RX�e��$X�,�������������_^��k��%M���wl��p��\�|W�
�ϟ�ٳgq��)ř3gp��i�8qǏW=z�V�2��~�?b߁8��aŁ#?�=?b���������.�-����މ�wm�7�v���
�Лw2ݱ_o�[vl�w�w�;�c��c�N�ر[�n�W_}�M_�/�l��l����|��[���X��[|�a�Y����e��j)�X�9�c�ֱd-o_�X��Ȣ5+���ԂU�2�g�5oӗ.D����<2w�LG�l��g�y�L�3��t�0�hjFiS�@TL���l���3��S�I��9oa SI*�TL#L+I)��)�P�D��P�<�Sڐ[߂���i��Z$�D)�_�&�T6#��IN�hAJU�;�V�!���IM+2j�� �)jY�ri�7�f2kg#�~.r�#�q>��[Uߦ�EM�)���I��*�GԤ:�!�b�]�М2g��/uҊ8\���`���Z���%�I�����R��"��!0CG��� ��C��I�U�_R�0� �(|X�P�tLԢ��C?7~��/=��gr_2
��ܯ�·p���@�Pۦ 0��PO��y�7/"�D�R�5P(<E�f�E<y<�'������mO$>�<GL�S
�||x>}��W�'�4�7��{��G������l�^�%ϸ��� ��$bS����d�#>��+�/��܆gJ>�����p8���	��Hȃgb>�(�^ܖ��7�ٛ���}���*�#r�(�!9�l��;���zd}�^�x�63U����lC9Ά��H��x���Mr�L��8��{�$L��,��9����ey��q<f��	�C{^����s�P����G�W<���'�:����s�����n�pM�W���p���ׅ�r�9v������l����I�2a���l8�x�yl�<N�$�G�MR�3�L�y��Mr���<X�X%�RN�`�uȸeB�5f�eGN�M.�X^O�:�&cbY#<
k��[�`��ǈ��9:x�K:�ϓ)���d�%TG
�4Qs�b �� "��������2��͘��"	"E���kI)��^>�Zk�P�lE�x�0��Q�4TÊ��%KN� �50l��QD�&NLR8N!7K�Qbn��Y)�k�Mz#��U�s���M�2��Q�[p_th�׮G3�:.�]&�O��4�zԼd9Ͳ�}�2�r��9P�d��դ���{J�C�0�O��ܩp$���\��)ϩ���v5�x�(Jj� ݎ����Mr�`�`�.�ד��7�~Ҕp�
16�A�7����s�"���)p�k������f��[<�[�E��*&N���>�:��E��W,�L�BP�lW�E��s]5��GX��M&5^����ݸ�M�E$bZV(⦭B��U�'�Nn���+�޺mˑE�ۖ���i[�ܶ��m]���(����b��՘�d����_V,�{,'+(�+мh>j��fM�L��z�l�-Z���K�B�n�M]�9�S�W}�v�܋�'/����=|��!�!=q�R;$�(�"�
��(�\���+����⟉���������W^iy�;�V;���eݺdǤ���;݁	#�~�|rp2__?�M�2����i]}}�WU�ϴt���io��t�����#t�Yo7:��v�3tr�O�Kd�\W����\C��-���~�������z��Ao�J�ww�޳����w�>�S>k�s:����4<�>>�~���������q��}\{|W��Շw�p��m\�w������7p��u��q��\��s�pH���Wq��5��qgo�ƹ�wp��=\���Ϲ��<�减q��n�)�=i����kO�"�ugn���[wq��}�É+�p��U:s��\Q道����%�;v��E�_��S�p��e9wU��tV���e���s8p�,�=��'�(��8�=GO��#'���S�{��Op��p����t�Z����{���g���3�9�m{bˏ��>lٳ����|�#�޽����������!�{�����u�D8m�Ar���6�������ZV����}D����]��ỽX�s֒/��L[�q�[6lf�%|C�ƲM��������W�k�}�F��^��;o�s_q[�|�u[��Za�������=VIe�[w�-Z�݅��`��o�T˒��2�'��`ɦo��o���-X�yV��7oŚo�q=;�n�Nl������bP��ܟ�d����Z�y���;��z'>�j�;��r+Vlྫྷ��Ȳ���?�`	�ɒ�_a��/1���X�v=���,�����ٲS÷;�z�woX�i+�<��l��o��Kn����j�s��|,����V�g�sW}��,Pf��3�����+0m�r�ԥ�вx)�?[��E���
L]�
Ӗ~��e�1M;<��\��6���6�ވ�ū0c)��k�0GX�Ż,դ���ƌϸ���fq��E+0e���^���P9]�ݹ�h���vʧ�A)m���N���ًQ;��]������u5.X�ƅK1y�|TΘ�ʙ\�̤|�,-�Q�܊¦6����(hlC�
��!��U��ܺ�H��WAt
h	�S9�Z�!������(@@J6����9����II/@Pj>�) �Ƞɟb�����`���?�*0+f�Ġ/�0�H��a��"=�$7N��T�	)�A�{�\�;�횜��'J�s"�n�))�0 I�'E�G.���P)qd ����c�7�B�$R����vW�n9Upe �� �fkS5\�x�w������`ܙ��lW�E�M�E�in��]������Vc��7D�e��<�Z&w2���ʖqY����`tR�5L,l�O��o��Y��4m,k��|ʚ�]��	^%M�,���e���*�!����چ^5C�%�z&����������ي��sG�k澥v#�%��CB�|$��GR��ܰɍd�"$7}���������K�ӖRv�!��+d�X�Ȟ�J�;k�f�D��/P�p�H����s���D��(��%�>C%����дt��%�Ѵ�|6S�1m�b��Z���d���1{�X�i#>��5fn�7oº�߱<܇�,��~���^v�+��
�A"�0��@�^Z	~5L�U�ƫ/)�#�c':t���~��w���ɰ��;�GC����������Ӄ��N<{���<A^�t���,/�,ߦ֡Ĕ2�CI�^���	/�ϰ�!����a�04�^
�f��~��Y$���w���o��n�<��!C�p����o�`��_0��k��
�:�wΧ�ٷ�s=�,�V��2���9����z^�{���st��1�u��~s�T�s?�ut�X��uK ���������_^�9�� ��?c��� �	�\���k��s/i�����w�w������5���z����y	�W0:�;���x����=�+A�Ч��^}�f����|��a`�ǩE����08���2� ����04	�4��0�!�=1�{���s�2�Z7��a���9��Z7��N8��zd�6d����,�e��k����hS�_���s�jY�����d	��X��g�G;�O�r=��u}�����[C7�<��SIOeߞw3P��t1���l[�-�DΟl���[wO/���`�Ӻ�65ە���y\o��u�}#�r�>��|n��'�ܟ'�O����HQ��}�%}�y�����s������O/���얼��Al'ק��K�V߯���Q��qu1Е ����=�π�	:�s�C��ץ��G�����{xn�y��9��缝练�39nIe�C��1��k��}y�� ��	ӧ�GO���c�:�~����~ro2�!�?�=�����{�<���綫S���΃�\{;�tt�k ���x�sN�I��Н/^�v����e����������t��}�xpOq�\�� �.�sW�e�#�z�.繏������>n����[��@�*�+7����+�|�-._��_Ź��q���9wg�_¹�2|���c'p��<�3�1��q��|��o+��[���m;�m�.l߹�?E��ꛭ�����k8���J3+W�ÊU바A�gK��3$���m�u�RL���3P�0��m(!��}2��_ӂ���ȫmF~}3
Ȥ�&55kh�
i�h��IM�0i�4\�a*��!�q�9-s�T$V�#a����ZD�V�!��!�%*(�n&f��+=�9j�'+�ٔ}��7I�� ���%\WY%"˫U^��Ɉ��U�����i�ejِ�RE0�A7웝��t�%�q_�F���}��"�_���r
�#��y��A��<�
T�*-�d2��8�4۫$U�^%�p>����4�E5*�EpqBJ�Vր@N��e]$dR�
jQX����D7(��4D7"����SqeM�@b�4d��"��� �AV�^��i�7���mY������
�/V�3�%o( ����p�2͢�2-���s��a�zԯXG֢�Ԯ�5+֠v��}��_�E�ڵhY�`y�j��֯@��嘾vf|!P|�R�W���5��`�:,��K,ذ�6n��o���m�b���n�9y'._�M�#�=�x������0�R;�R��u���%y+�#��#���Q�u�<�����t���H�c�����5��ye� �DTRc��%��Y���X}�D��H�s��5��J�ϓ��8�t]��Y��&�m�v�|��WBƂ����R�iRhK�H�� T��U��H���`!����Я��;h��q
j����V�I7�L
p�������2��ZV���UM7@j��(Z}�j������K����t�����KI�H�q���/�����I�x�Dzu������Oz��_=�N/�K�?%��b�ǂ���E����]O������g��� ��t��d   IDATqX�;��E��x�T�9_�c��=��oy��i�S��D�I	�y���@�3>:04Ё�~aP6�����y�(8
��f�Ϟ�x��x��y�{I������l���ӻxQ�8���]�����A$R�H���m	��n^_���v޳�n�S�c�<��?��5�upC\~�����%��
�s
i��NZe;�I��٫�G]�6D�i��}U�s�s�F�짘?����g���|�Z^I_2�x��xI^?��A��W~��^�@7���ޗ2�K/y�	����V/�9܏���A�P��7r_��0��c��������k"�N�u�y�~�x5�<M�:޿��;;�r�\'�=H�x�j��m���W����z���6y�zx��\gm�-�כ B�?D��A�˰3y�=�|��q>��|��	�����CD=���l��}�9���z��c��w������MD�&�</~V����y�K�����|��*�	�a�×��/��� ���=��C��\�.ޓ�L��G��ȼ�Tk���̫YN�l'�U7�>�����aM^ǀ������T�)�tY���Vx��i�L��6�<�?g?�*�8�dk��/�r�u�ؒc���J�lR�c[�lK��D]93���� ����}~��H��I����o7�o�9¹ލ�8 }��n6qP�#�6z][�߮݃�{vucî��W��v���M�r��}��n��s�n��n�o���p��uw-.ݸF�k�յ��/�^�/��x�.\[����y�ϯ_����|µ磯/��}j�>�������7�������A�m�?�{������:~�<�ĥ��������������/\��߼n�o\�O)��+��/����9̟.~����W�����ěg��_�c���Ͻv�^:�?+θ8/�欝|�7���o�/V�V�|g͡sw����7�؋����������rZ�u</{�#���ճ���e?��y����c}���O���??a����{�^�;�����_�3/��?:�/ �������g�ߒgu�D�<���<m?��|�o���P�g�?uR�?���Ͽb�?���๓�{���T?P=��;-~t��%Ͻ�[{^�]�����ى5x�];q�=;/�����|�~�Ư���u�|�{��6>wƎ�K��Kۼ���z�v�S�"���h�sv����ڟpD�b}�.ܢ_oܶ[[�A��x��.�[������:
W�i-�8��ta3��To��Z��9hVt����a�/�Wȋa/z��j���M;����Py:b�9i��6��ك
&�5#F�kFh��Λc�����aO[,�hUy$�����8q�<)���SJ�R�T	��BR�����D �	�A�:/��aR�f0���6����ψ��pfrC0��~�O�Q=�%�Y�IBȓ3	:���_Zy�49ΕV�T:�+J!b#���Ĥ�2Uv�X�p*2D��o�3K�8EB<��Հ�$�<FL:���8Gp��9Jv,���vS����L�S&���L�5hC
�KوV�b�DTN����O`��2���'���`Dq�HO�I�!/~��P}�s@D>L�Ϙ!�3�d� �6��t 0�#�e_����	�r�E#�Ӥ���F�}�\�cҗ�SN�p�(��Q��K�iE[m����.�@XxJ�ҏ�^8QN�R_�)�NBu!�(eO�`�HEJ��6řȱiN{��Di�(-�c��a^"X爘�4G1Ch5"�gCh�c�)�K87������,P��\`��� W����;�v:�&�	ol��~	uW�1�Vb�R��s��Q)(�"LLȻ"oDzF�G&������#�d�S�s�>�$E�g�>���Ʋ�%dO9`j?�W��A���;�� ���g��9 �N���υ·��RF$�22�J.D������8e	Ϙ�!���';�-�q�R9�@����-��;��p��=�4l����C� ���{�>}lѧN"R�����bb�����j%��6�α�1�['�%�SKqPt�t�3�6C�cH�h�d�h�!��s�|J�y� �A�ݢ��-�c��̤�����h��4�q��^�{TП�䔌Sケ�-�0��ˎ[�h���r"xtԵ���)h���q<�sNNH���X���RJ�v}��]���-ڰ�E�m C������B��W(���g������1�O "�3}hXO�C��3\��3��%ۻC{�����C�"M�<zQ�bsǧ�c���<Ǯ=���1i=�\o������|�0�%o�I�]��}���tmc�cwo��G�����v��=�;v囻�܁�����?|d7mڍMxL���e��ɣӱ[u}��o8�����,�o�c�w�v��mWi��7����v��7���;�������;8Ew��������M�x�]�w�.m�@�^�+�o���)�=���>&�浞�i��J�ﷅ�a1,!��3D0��{�>D,��3#�כm�Z���CZU:Vz���Gq�0qTeW���G=���)��=�.TȞ���k�d���ټ��c�ÌYB��!��P����^��-A�E���y���g/F�֪s]V6E��|%H)��!�8sT�OR:��;z�3ҵ�X.��b%��'/������{��3X	i�=�nSD{�`�W�4�74�X��'�W!�ʦ�[0���*���S,��3f#ʱ�0,�E�;R��S~�ӹV�"��ɠ�Lz���C&pM�Q�M&�4���Ѭ��pqc�iE��	&�T>"Bu��V������7��	�ӥ��)�G�xx.ʎq�������`�d�@�y1 ��~�a*�(4YP���Bʍ��`V�N�����]eO�ٗ�0�4���B廭�t�|��/Z��W��c�oPO�Y{޻�]�v�Q�/qE{�8�|7u����iӐr��Ǡ��?\m��6�E��0�(O���đDOBl�0����Yi�V[�S����%�]�U"��<�R� P�MB_��WP�#ZDF��4)�F[3�%#��ޝ�w*�y�"�Eg��rK����k�}��Be��:i���*A ���MB�%`�0�V���v��{���!m4�-���>���2�Y��-`�������cHX�Q[Gl���p_��i�;^MGk�ϒ�C����!��6	b��g�,h;Ւ<����/�u)a|Y��S���h�x
5�6���O�I��]�	�W���0�����H���  �9���s���	ϣ�Oѳ��vI��� ���M�;]����v��{ѱ�so��`�X���~����h��v
�u#�Rl���#����e]��/�q>�9�<����U\W�Gs��! ��i~�ܜ�4�O�Ii�����C�9ut�#�m#8SD���q36s �m�����͊���ġ�����gě+�i�����V���唹qΜ�`��c�{��@P��a�'�Dl�3�����j}y�|�9bN�boZ�h��@MN��a�Mh�BmM�@�p]뫒���r�8�'�%����K��.�����j�p>��+q�Ę�*����7tԭ�����x*+������2r�3ҥ�i��XN�#�����g�|�*�f(3��E��V{�/(w�SՈ���f
+���ۃ}����#N���m�����J�2?�"^�E������h�b&�)q*1� �"P�9'�9�Q[,�HXJj�X�+j΅˗<��o���Jhkcʀ��3~�`�=ő v[-xG
�V	a��JغŽ�ŷ^��^5m�K��/_�� H3��3�A�j�x��9H�X��<�eJ�j�Z3hO�T%�+<�	YH?%>�>q�S7��V�ܪ�R�rM\�u��O�­�铬D0�	e���k�	�C���K�%4�̈́�L��#��"��f{
�����)����vi��A�0!��S�=���!�R`j�h�C\�V�_(MN[d��(1�ں�V<t
��0��?b�DL߈hߐ��'�?������{bH��D	��.C�ѤҦ�Ĵq���p�=���Ct$ψ�"���=
�Ő�����g"�&;*AX�?]{�%��x�P"l���N䔙��;�`��TaG���<�G�,���)���k���Y$U��^{������#a�l����:�jٞp�kg+��ϲ_�-d=sB�Ŵ�������C���Ő�	��U�2�	oG����k�U�ĐpO��q�kH�\��� ��6V]��U~��(á~����H��1���*�:����^�/@u��V�y�ae�x�3�:j+R-$0��0ΰŀ�ɐ�8`L��Ҋ��?�\�qƄO�*�A�L�IE9�a(�%T.�;Q>�%��䈶fGt��Os@�ݴJ���e�8����A�q���1��8�q�� ��>)�L{k+Hθ�� i�s+���]�ێ�y�ti$��#B7DXB0�BuӸ0+R�}֨�	vZ��nc��� ��#ZW4acl��L�GNPG�c���P��`��P�{�i<ZQG�O�*��T�����!�w�zCǔ:4��8�9�f��s�2��M�������9S��c͜�f���h�=�ςwsFLi���5cws��	-F�G6�Q�D6ׂ����0mA�ס07���s�a�E�/:�Z_�6��GX�̓.�/@	-NU���+�('ާ���Xη..�q���I_S}��9��q�8�L"݆x]� �bY�&8��
�.��s������(�x�$�qjt���'�4��(��S��m1��J�.�Ä���A�·M�k��� GA�u)�    IEND�B`�PK    S�U��V��       jsons/user_defined.json���n�0E%��D��(�x�EӢ�UaE�Q������0~!���Q�9spgt��hXu�����2�mM�f��u-\�I�8��2��h�c��W�������fa��Q+(�j0ί�}��bG^ΐ���ʕ %�I.��s�פ`E)U�'�ڷ�?����鵷ݰy����H|ҵ��������Q;>�F�u�(;�}qO��� �k[�{	�]�u����P�z�~����&���a�%��"�"�h�/�}?k�J:�fvN.��8�U����%:9'=��]��җ����5��`�y�?�g��i�^� ���?u���k��|��S�*QaZ0���:�8��	י�z��c��<�'�m���x�g,!��ٻ9�Ȇ�O�'<{:9�|����l�v��.��گ�O��^��ց̈ܔENeY@0՘�Y��U8�V��ε6r����nէbCҤ�`���!��I���rs�����PK
    S�U&!S  �                   cirkitFile.jsonPK
   �jgUD�#��9 �9 /             �  images/44ae2a6d-294a-417e-8c08-7c32f15c3a8c.pngPK
   �kgU�g<��4 v; /             �K images/b9728b98-ae2c-4f30-943d-a61b81bf7cce.pngPK
   @jgU�\���	 2	 /             ƀ images/ee25a61b-6355-4858-a778-65c1949b8af0.pngPK
    S�U��V��                 � jsons/user_defined.jsonPK      �  �   